<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-124.657,32.6416,219.936,-143.531</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>54.5,-4.5</position>
<gparam>LABEL_TEXT Front Panel</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AI_XOR4</type>
<position>19,-18.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>128 </input>
<input>
<ID>IN_2</ID>251 </input>
<input>
<ID>IN_3</ID>250 </input>
<output>
<ID>OUT</ID>740 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>7.5,-12</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>1,-24.5</position>
<output>
<ID>OUT_0</ID>250 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>DE_TO</type>
<position>39,-18.5</position>
<input>
<ID>IN_0</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>264</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>71,-33</position>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>273 </input>
<input>
<ID>IN_2</ID>274 </input>
<input>
<ID>IN_3</ID>275 </input>
<input>
<ID>IN_4</ID>276 </input>
<input>
<ID>IN_5</ID>277 </input>
<input>
<ID>IN_6</ID>278 </input>
<input>
<ID>IN_7</ID>279 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 223</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>266</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>117.5,-31</position>
<input>
<ID>IN_0</ID>263 </input>
<input>
<ID>IN_1</ID>264 </input>
<input>
<ID>IN_2</ID>266 </input>
<input>
<ID>IN_3</ID>267 </input>
<input>
<ID>IN_4</ID>268 </input>
<input>
<ID>IN_5</ID>269 </input>
<input>
<ID>IN_6</ID>270 </input>
<input>
<ID>IN_7</ID>271 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>268</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>108,-59.5</position>
<input>
<ID>IN_0</ID>312 </input>
<input>
<ID>IN_1</ID>286 </input>
<input>
<ID>IN_2</ID>285 </input>
<input>
<ID>IN_3</ID>284 </input>
<input>
<ID>IN_4</ID>283 </input>
<input>
<ID>IN_5</ID>282 </input>
<input>
<ID>IN_6</ID>281 </input>
<input>
<ID>IN_7</ID>280 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>270</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>67,-63</position>
<input>
<ID>IN_0</ID>330 </input>
<input>
<ID>IN_1</ID>316 </input>
<input>
<ID>IN_2</ID>314 </input>
<input>
<ID>IN_3</ID>313 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>272</ID>
<type>AA_TOGGLE</type>
<position>1.5,-52</position>
<output>
<ID>OUT_0</ID>248 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>274</ID>
<type>DE_TO</type>
<position>13.5,-52</position>
<input>
<ID>IN_0</ID>248 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>662</ID>
<type>GA_LED</type>
<position>107.5,-8</position>
<input>
<ID>N_in0</ID>720 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>278</ID>
<type>DA_FROM</type>
<position>2,-20.5</position>
<input>
<ID>IN_0</ID>251 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck3</lparam></gate>
<gate>
<ID>670</ID>
<type>DA_FROM</type>
<position>104,-8</position>
<input>
<ID>IN_0</ID>720 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>672</ID>
<type>GA_LED</type>
<position>107.5,-12</position>
<input>
<ID>N_in0</ID>721 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>674</ID>
<type>DA_FROM</type>
<position>104,-12</position>
<input>
<ID>IN_0</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Execute</lparam></gate>
<gate>
<ID>294</ID>
<type>DA_FROM</type>
<position>47.5,-22</position>
<input>
<ID>IN_0</ID>279 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>295</ID>
<type>DA_FROM</type>
<position>48,-25.5</position>
<input>
<ID>IN_0</ID>278 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>296</ID>
<type>DA_FROM</type>
<position>48,-28</position>
<input>
<ID>IN_0</ID>277 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>297</ID>
<type>DA_FROM</type>
<position>49,-31</position>
<input>
<ID>IN_0</ID>276 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>298</ID>
<type>DA_FROM</type>
<position>50,-34</position>
<input>
<ID>IN_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>299</ID>
<type>DA_FROM</type>
<position>49,-36.5</position>
<input>
<ID>IN_0</ID>274 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>300</ID>
<type>DA_FROM</type>
<position>47,-39.5</position>
<input>
<ID>IN_0</ID>273 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>301</ID>
<type>DA_FROM</type>
<position>47,-43</position>
<input>
<ID>IN_0</ID>272 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>302</ID>
<type>DA_FROM</type>
<position>96.5,-16.5</position>
<input>
<ID>IN_0</ID>271 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>303</ID>
<type>DA_FROM</type>
<position>96.5,-20</position>
<input>
<ID>IN_0</ID>270 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>304</ID>
<type>DA_FROM</type>
<position>97,-22.5</position>
<input>
<ID>IN_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>305</ID>
<type>DA_FROM</type>
<position>97,-25.5</position>
<input>
<ID>IN_0</ID>268 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>306</ID>
<type>DA_FROM</type>
<position>97,-28.5</position>
<input>
<ID>IN_0</ID>267 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>307</ID>
<type>DA_FROM</type>
<position>97,-31</position>
<input>
<ID>IN_0</ID>266 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>308</ID>
<type>DA_FROM</type>
<position>96.5,-34.5</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>309</ID>
<type>DA_FROM</type>
<position>97,-38</position>
<input>
<ID>IN_0</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>312</ID>
<type>DA_FROM</type>
<position>55,-57</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 11</lparam></gate>
<gate>
<ID>313</ID>
<type>DA_FROM</type>
<position>53,-62</position>
<input>
<ID>IN_0</ID>314 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 10</lparam></gate>
<gate>
<ID>314</ID>
<type>DA_FROM</type>
<position>52,-65.5</position>
<input>
<ID>IN_0</ID>316 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 9</lparam></gate>
<gate>
<ID>315</ID>
<type>DA_FROM</type>
<position>51.5,-69</position>
<input>
<ID>IN_0</ID>330 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 8</lparam></gate>
<gate>
<ID>316</ID>
<type>DA_FROM</type>
<position>93.5,-48.5</position>
<input>
<ID>IN_0</ID>280 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 7</lparam></gate>
<gate>
<ID>317</ID>
<type>DA_FROM</type>
<position>94,-54</position>
<input>
<ID>IN_0</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 6</lparam></gate>
<gate>
<ID>318</ID>
<type>DA_FROM</type>
<position>94.5,-57</position>
<input>
<ID>IN_0</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 5</lparam></gate>
<gate>
<ID>319</ID>
<type>DA_FROM</type>
<position>95,-59.5</position>
<input>
<ID>IN_0</ID>283 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 4</lparam></gate>
<gate>
<ID>320</ID>
<type>DA_FROM</type>
<position>94.5,-61.5</position>
<input>
<ID>IN_0</ID>284 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 3</lparam></gate>
<gate>
<ID>321</ID>
<type>DA_FROM</type>
<position>95.5,-65</position>
<input>
<ID>IN_0</ID>285 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 2</lparam></gate>
<gate>
<ID>322</ID>
<type>DA_FROM</type>
<position>96,-68</position>
<input>
<ID>IN_0</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 1</lparam></gate>
<gate>
<ID>323</ID>
<type>DA_FROM</type>
<position>95,-72.5</position>
<input>
<ID>IN_0</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 0</lparam></gate>
<gate>
<ID>148</ID>
<type>DA_FROM</type>
<position>6,-17.5</position>
<input>
<ID>IN_0</ID>128 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck2</lparam></gate>
<gate>
<ID>746</ID>
<type>BB_CLOCK</type>
<position>5,-29.5</position>
<output>
<ID>CLK</ID>742 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 25</lparam></gate>
<gate>
<ID>753</ID>
<type>AI_XOR2</type>
<position>30.5,-22.5</position>
<input>
<ID>IN_0</ID>740 </input>
<input>
<ID>IN_1</ID>741 </input>
<output>
<ID>OUT</ID>739 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>755</ID>
<type>AA_AND2</type>
<position>19,-30.5</position>
<input>
<ID>IN_0</ID>742 </input>
<input>
<ID>IN_1</ID>743 </input>
<output>
<ID>OUT</ID>741 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>757</ID>
<type>AA_TOGGLE</type>
<position>6.5,-36.5</position>
<output>
<ID>OUT_0</ID>743 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>759</ID>
<type>AA_LABEL</type>
<position>1,-36</position>
<gparam>LABEL_TEXT Run</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9.5,-12,16,-12</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>16 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>16,-15.5,16,-12</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-52,11.5,-52</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<connection>
<GID>272</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-24.5,11.5,-21.5</points>
<intersection>-24.5 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-21.5,16,-21.5</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3,-24.5,11.5,-24.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-20.5,16,-20.5</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>16 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,-20.5,16,-19.5</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>-20.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,-38,109,-34</points>
<intersection>-38 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109,-34,112.5,-34</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-38,109,-38</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>109 0</intersection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-34.5,107,-33</points>
<intersection>-34.5 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-33,112.5,-33</points>
<connection>
<GID>266</GID>
<name>IN_1</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98.5,-34.5,107,-34.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-32,107,-31</points>
<intersection>-32 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-32,112.5,-32</points>
<connection>
<GID>266</GID>
<name>IN_2</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-31,107,-31</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-31,107.5,-28.5</points>
<intersection>-31 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-31,112.5,-31</points>
<connection>
<GID>266</GID>
<name>IN_3</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-28.5,107.5,-28.5</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-30,108.5,-25.5</points>
<intersection>-30 1</intersection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-30,112.5,-30</points>
<connection>
<GID>266</GID>
<name>IN_4</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-25.5,108.5,-25.5</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-29,109.5,-22.5</points>
<intersection>-29 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-29,112.5,-29</points>
<connection>
<GID>266</GID>
<name>IN_5</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-22.5,109.5,-22.5</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-28,110,-20</points>
<intersection>-28 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-28,112.5,-28</points>
<connection>
<GID>266</GID>
<name>IN_6</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98.5,-20,110,-20</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-27,111.5,-16.5</points>
<intersection>-27 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,-27,112.5,-27</points>
<connection>
<GID>266</GID>
<name>IN_7</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98.5,-16.5,111.5,-16.5</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-43,63,-36</points>
<intersection>-43 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-36,66,-36</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-43,63,-43</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-39.5,61,-35</points>
<intersection>-39.5 2</intersection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-35,66,-35</points>
<connection>
<GID>264</GID>
<name>IN_1</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-39.5,61,-39.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-36.5,60,-34</points>
<intersection>-36.5 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60,-34,66,-34</points>
<connection>
<GID>264</GID>
<name>IN_2</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-36.5,60,-36.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-34,58,-33</points>
<intersection>-34 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-33,66,-33</points>
<connection>
<GID>264</GID>
<name>IN_3</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-34,58,-34</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-32,58,-31</points>
<intersection>-32 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-32,66,-32</points>
<connection>
<GID>264</GID>
<name>IN_4</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-31,58,-31</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-31,60.5,-28</points>
<intersection>-31 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-31,66,-31</points>
<connection>
<GID>264</GID>
<name>IN_5</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-28,60.5,-28</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-30,61,-25.5</points>
<intersection>-30 1</intersection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-30,66,-30</points>
<connection>
<GID>264</GID>
<name>IN_6</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-25.5,61,-25.5</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-29,62,-22</points>
<intersection>-29 1</intersection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-29,66,-29</points>
<connection>
<GID>264</GID>
<name>IN_7</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-22,62,-22</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-55.5,102,-48.5</points>
<intersection>-55.5 1</intersection>
<intersection>-48.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-55.5,103,-55.5</points>
<connection>
<GID>268</GID>
<name>IN_7</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,-48.5,102,-48.5</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-56.5,101,-54</points>
<intersection>-56.5 1</intersection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-56.5,103,-56.5</points>
<connection>
<GID>268</GID>
<name>IN_6</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96,-54,101,-54</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96.5,-57,103,-57</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>103 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>103,-57.5,103,-57</points>
<connection>
<GID>268</GID>
<name>IN_5</name></connection>
<intersection>-57 1</intersection></vsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-59.5,101,-58.5</points>
<intersection>-59.5 2</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-58.5,103,-58.5</points>
<connection>
<GID>268</GID>
<name>IN_4</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-59.5,101,-59.5</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-61.5,100,-59.5</points>
<intersection>-61.5 2</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-59.5,103,-59.5</points>
<connection>
<GID>268</GID>
<name>IN_3</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-61.5,100,-61.5</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-65,100.5,-60.5</points>
<intersection>-65 2</intersection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-60.5,103,-60.5</points>
<connection>
<GID>268</GID>
<name>IN_2</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-65,100.5,-65</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-68,101,-61.5</points>
<intersection>-68 2</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-61.5,103,-61.5</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98,-68,101,-68</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-72.5,102,-62.5</points>
<intersection>-72.5 2</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-62.5,103,-62.5</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-72.5,102,-72.5</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-61,60.5,-57</points>
<intersection>-61 1</intersection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-61,64,-61</points>
<connection>
<GID>270</GID>
<name>IN_3</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-57,60.5,-57</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-62,64,-62</points>
<connection>
<GID>270</GID>
<name>IN_2</name></connection>
<connection>
<GID>313</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-65.5,60.5,-63</points>
<intersection>-65.5 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-63,64,-63</points>
<connection>
<GID>270</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-65.5,60.5,-65.5</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8,-17.5,16,-17.5</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>16 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>16,-17.5,16,-17.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-69,61,-64</points>
<intersection>-69 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-64,64,-64</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-69,61,-69</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>720</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106,-8,106.5,-8</points>
<connection>
<GID>662</GID>
<name>N_in0</name></connection>
<connection>
<GID>670</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>721</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106,-12,106.5,-12</points>
<connection>
<GID>672</GID>
<name>N_in0</name></connection>
<connection>
<GID>674</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>739</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-22.5,35,-18.5</points>
<intersection>-22.5 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-18.5,37,-18.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-22.5,35,-22.5</points>
<connection>
<GID>753</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>740</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-21.5,25,-18.5</points>
<intersection>-21.5 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-21.5,27.5,-21.5</points>
<connection>
<GID>753</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-18.5,25,-18.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>741</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-30.5,24.5,-23.5</points>
<intersection>-30.5 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-23.5,27.5,-23.5</points>
<connection>
<GID>753</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-30.5,24.5,-30.5</points>
<connection>
<GID>755</GID>
<name>OUT</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>742</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9,-29.5,16,-29.5</points>
<connection>
<GID>755</GID>
<name>IN_0</name></connection>
<connection>
<GID>746</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>743</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-36.5,12,-31.5</points>
<intersection>-36.5 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-31.5,16,-31.5</points>
<connection>
<GID>755</GID>
<name>IN_1</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-36.5,12,-36.5</points>
<connection>
<GID>757</GID>
<name>OUT_0</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-44.7154,9.28712,192.619,-112.05</PageViewport>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>57.5,6.5</position>
<gparam>LABEL_TEXT Memory</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AI_RAM_12x16</type>
<position>55,-27</position>
<input>
<ID>ADDRESS_0</ID>19 </input>
<input>
<ID>ADDRESS_1</ID>18 </input>
<input>
<ID>ADDRESS_10</ID>9 </input>
<input>
<ID>ADDRESS_11</ID>8 </input>
<input>
<ID>ADDRESS_2</ID>17 </input>
<input>
<ID>ADDRESS_3</ID>16 </input>
<input>
<ID>ADDRESS_4</ID>15 </input>
<input>
<ID>ADDRESS_5</ID>14 </input>
<input>
<ID>ADDRESS_6</ID>13 </input>
<input>
<ID>ADDRESS_7</ID>12 </input>
<input>
<ID>ADDRESS_8</ID>11 </input>
<input>
<ID>ADDRESS_9</ID>10 </input>
<input>
<ID>DATA_IN_0</ID>28 </input>
<input>
<ID>DATA_IN_1</ID>29 </input>
<input>
<ID>DATA_IN_10</ID>25 </input>
<input>
<ID>DATA_IN_11</ID>24 </input>
<input>
<ID>DATA_IN_12</ID>23 </input>
<input>
<ID>DATA_IN_13</ID>22 </input>
<input>
<ID>DATA_IN_14</ID>21 </input>
<input>
<ID>DATA_IN_15</ID>20 </input>
<input>
<ID>DATA_IN_2</ID>30 </input>
<input>
<ID>DATA_IN_3</ID>31 </input>
<input>
<ID>DATA_IN_4</ID>32 </input>
<input>
<ID>DATA_IN_5</ID>33 </input>
<input>
<ID>DATA_IN_6</ID>34 </input>
<input>
<ID>DATA_IN_7</ID>35 </input>
<input>
<ID>DATA_IN_8</ID>27 </input>
<input>
<ID>DATA_IN_9</ID>26 </input>
<output>
<ID>DATA_OUT_0</ID>28 </output>
<output>
<ID>DATA_OUT_1</ID>29 </output>
<output>
<ID>DATA_OUT_10</ID>25 </output>
<output>
<ID>DATA_OUT_11</ID>24 </output>
<output>
<ID>DATA_OUT_12</ID>23 </output>
<output>
<ID>DATA_OUT_13</ID>22 </output>
<output>
<ID>DATA_OUT_14</ID>21 </output>
<output>
<ID>DATA_OUT_15</ID>20 </output>
<output>
<ID>DATA_OUT_2</ID>30 </output>
<output>
<ID>DATA_OUT_3</ID>31 </output>
<output>
<ID>DATA_OUT_4</ID>32 </output>
<output>
<ID>DATA_OUT_5</ID>33 </output>
<output>
<ID>DATA_OUT_6</ID>34 </output>
<output>
<ID>DATA_OUT_7</ID>35 </output>
<output>
<ID>DATA_OUT_8</ID>27 </output>
<output>
<ID>DATA_OUT_9</ID>26 </output>
<input>
<ID>ENABLE_0</ID>7 </input>
<input>
<ID>write_clock</ID>1 </input>
<input>
<ID>write_enable</ID>6 </input>
<gparam>angle 0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:0 49156</lparam>
<lparam>Address:1 57343</lparam>
<lparam>Address:2 65022</lparam>
<lparam>Address:3 57344</lparam></gate>
<gate>
<ID>8</ID>
<type>DA_FROM</type>
<position>88,-22</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>22</ID>
<type>DA_FROM</type>
<position>82,-26.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Mem Write</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>83.5,-31</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Mem Read</lparam></gate>
<gate>
<ID>26</ID>
<type>DA_FROM</type>
<position>30,-7.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 11</lparam></gate>
<gate>
<ID>27</ID>
<type>DA_FROM</type>
<position>30,-10.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 10</lparam></gate>
<gate>
<ID>28</ID>
<type>DA_FROM</type>
<position>28.5,-13.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 9</lparam></gate>
<gate>
<ID>29</ID>
<type>DA_FROM</type>
<position>28.5,-17</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 8</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>28.5,-19.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 7</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>28.5,-22</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 6</lparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>29.5,-24.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 5</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>29,-27</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 4</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>29.5,-29.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 3</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>29.5,-32</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 2</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>29.5,-35</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 1</lparam></gate>
<gate>
<ID>37</ID>
<type>DA_FROM</type>
<position>29.5,-37.5</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Addr 0</lparam></gate>
<gate>
<ID>39</ID>
<type>DE_TO</type>
<position>29.5,-41.5</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>29.5,-44.5</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>41</ID>
<type>DE_TO</type>
<position>29,-47.5</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>29,-51</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>43</ID>
<type>DE_TO</type>
<position>29,-54</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>28.5,-56.5</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_TO</type>
<position>27,-59.5</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>27.5,-64</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>73.5,-42</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>49</ID>
<type>DE_TO</type>
<position>73.5,-44.5</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>50</ID>
<type>DE_TO</type>
<position>73,-48</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>51</ID>
<type>DE_TO</type>
<position>73,-51</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>52</ID>
<type>DE_TO</type>
<position>73,-54</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>53</ID>
<type>DE_TO</type>
<position>72.5,-56.5</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>54</ID>
<type>DE_TO</type>
<position>73,-59</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>55</ID>
<type>DE_TO</type>
<position>73,-63</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,-22,86,-22</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>64 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>64,-25.5,64,-22</points>
<connection>
<GID>6</GID>
<name>write_clock</name></connection>
<intersection>-22 1</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,-26.5,80,-26.5</points>
<connection>
<GID>6</GID>
<name>write_enable</name></connection>
<connection>
<GID>22</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-31,68,-27.5</points>
<intersection>-31 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-27.5,68,-27.5</points>
<connection>
<GID>6</GID>
<name>ENABLE_0</name></connection>
<intersection>68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-31,81.5,-31</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-7.5,46,-7.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>46 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>46,-21.5,46,-7.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_11</name></connection>
<intersection>-7.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-22.5,45,-10.5</points>
<intersection>-22.5 1</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-22.5,46,-22.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_10</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-10.5,45,-10.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-23.5,44,-13.5</points>
<intersection>-23.5 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-23.5,46,-23.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_9</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-13.5,44,-13.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-17,43.5,-17</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>43.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43.5,-24.5,43.5,-17</points>
<intersection>-24.5 4</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>43.5,-24.5,46,-24.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_8</name></connection>
<intersection>43.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-25.5,40,-19.5</points>
<intersection>-25.5 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-25.5,46,-25.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_7</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-19.5,40,-19.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-26.5,46,-26.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_6</name></connection>
<intersection>38 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>38,-26.5,38,-22</points>
<intersection>-26.5 1</intersection>
<intersection>-22 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>30.5,-22,38,-22</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>38 3</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-27.5,37,-24.5</points>
<intersection>-27.5 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-27.5,46,-27.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_5</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-24.5,37,-24.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-28.5,35.5,-27</points>
<intersection>-28.5 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-28.5,46,-28.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_4</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-27,35.5,-27</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-29.5,46,-29.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_3</name></connection>
<connection>
<GID>34</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-32,41.5,-30.5</points>
<intersection>-32 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-30.5,46,-30.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_2</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-32,41.5,-32</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-35,43,-31.5</points>
<intersection>-35 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-31.5,46,-31.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_1</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-35,43,-35</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-37.5,45,-32.5</points>
<intersection>-37.5 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-32.5,46,-32.5</points>
<connection>
<GID>6</GID>
<name>ADDRESS_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-37.5,45,-37.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-41.5,47.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_15</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_15</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-41.5,47.5,-41.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-44.5,48.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_14</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_14</name></connection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-44.5,48.5,-44.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-47.5,49.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_13</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_13</name></connection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-47.5,49.5,-47.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-51,50.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_12</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_12</name></connection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-51,50.5,-51</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-54,51.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_11</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_11</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-54,51.5,-54</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-56.5,52.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_10</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_10</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-56.5,52.5,-56.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-59.5,53.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_9</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_9</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-59.5,53.5,-59.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-64,54.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_8</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_8</name></connection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-64,54.5,-64</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-42,62.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_0</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-42,71.5,-42</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-44.5,61.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_1</name></connection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-44.5,71.5,-44.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-48,60.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_2</name></connection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-48,71,-48</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-51,59.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_3</name></connection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-51,71,-51</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-54,58.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_4</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-54,71,-54</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-56.5,57.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_5</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-56.5,70.5,-56.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-59,56.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_6</name></connection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-59,71,-59</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-63,55.5,-38</points>
<connection>
<GID>6</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>6</GID>
<name>DATA_IN_7</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-63,71,-63</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-56.9158,19.5548,180.419,-101.782</PageViewport>
<gate>
<ID>772</ID>
<type>DE_TO</type>
<position>104.5,-68</position>
<input>
<ID>IN_0</ID>681 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I1</lparam></gate>
<gate>
<ID>773</ID>
<type>DE_TO</type>
<position>106.5,-68</position>
<input>
<ID>IN_0</ID>682 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I2</lparam></gate>
<gate>
<ID>774</ID>
<type>DE_TO</type>
<position>108.5,-68</position>
<input>
<ID>IN_0</ID>683 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I3</lparam></gate>
<gate>
<ID>775</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>114,-61</position>
<input>
<ID>ENABLE_0</ID>693 </input>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>70 </input>
<output>
<ID>OUT_0</ID>684 </output>
<output>
<ID>OUT_1</ID>685 </output>
<output>
<ID>OUT_2</ID>686 </output>
<output>
<ID>OUT_3</ID>687 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>776</ID>
<type>DE_TO</type>
<position>111.5,-68</position>
<input>
<ID>IN_0</ID>684 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I4</lparam></gate>
<gate>
<ID>777</ID>
<type>DE_TO</type>
<position>113.5,-68</position>
<input>
<ID>IN_0</ID>685 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I5</lparam></gate>
<gate>
<ID>778</ID>
<type>DE_TO</type>
<position>115.5,-68</position>
<input>
<ID>IN_0</ID>686 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I6</lparam></gate>
<gate>
<ID>779</ID>
<type>DE_TO</type>
<position>117.5,-68</position>
<input>
<ID>IN_0</ID>687 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I7</lparam></gate>
<gate>
<ID>780</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>129,-61</position>
<input>
<ID>ENABLE_0</ID>700 </input>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>65 </input>
<input>
<ID>IN_3</ID>66 </input>
<output>
<ID>OUT_0</ID>688 </output>
<output>
<ID>OUT_1</ID>689 </output>
<output>
<ID>OUT_2</ID>690 </output>
<output>
<ID>OUT_3</ID>691 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>781</ID>
<type>DE_TO</type>
<position>124,-73</position>
<input>
<ID>IN_0</ID>688 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I8</lparam></gate>
<gate>
<ID>782</ID>
<type>DE_TO</type>
<position>127,-73</position>
<input>
<ID>IN_0</ID>689 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I9</lparam></gate>
<gate>
<ID>783</ID>
<type>DE_TO</type>
<position>129.5,-72.5</position>
<input>
<ID>IN_0</ID>690 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I10</lparam></gate>
<gate>
<ID>784</ID>
<type>DE_TO</type>
<position>132,-73.5</position>
<input>
<ID>IN_0</ID>691 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I11</lparam></gate>
<gate>
<ID>785</ID>
<type>DA_FROM</type>
<position>119,-61</position>
<input>
<ID>IN_0</ID>693 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID IR-PC</lparam></gate>
<gate>
<ID>786</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>139.5,-70</position>
<input>
<ID>ENABLE_0</ID>699 </input>
<input>
<ID>IN_0</ID>698 </input>
<input>
<ID>IN_1</ID>698 </input>
<input>
<ID>IN_2</ID>698 </input>
<input>
<ID>IN_3</ID>698 </input>
<output>
<ID>OUT_0</ID>694 </output>
<output>
<ID>OUT_1</ID>695 </output>
<output>
<ID>OUT_2</ID>696 </output>
<output>
<ID>OUT_3</ID>697 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>787</ID>
<type>DE_TO</type>
<position>136,-82</position>
<input>
<ID>IN_0</ID>694 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I8</lparam></gate>
<gate>
<ID>788</ID>
<type>DE_TO</type>
<position>139,-81.5</position>
<input>
<ID>IN_0</ID>695 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I9</lparam></gate>
<gate>
<ID>789</ID>
<type>DE_TO</type>
<position>143.5,-81</position>
<input>
<ID>IN_0</ID>696 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I10</lparam></gate>
<gate>
<ID>790</ID>
<type>DE_TO</type>
<position>147,-81.5</position>
<input>
<ID>IN_0</ID>697 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I11</lparam></gate>
<gate>
<ID>792</ID>
<type>BA_TRI_STATE</type>
<position>140.5,-63</position>
<input>
<ID>ENABLE_0</ID>699 </input>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>698 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>793</ID>
<type>DA_FROM</type>
<position>150,-70</position>
<input>
<ID>IN_0</ID>699 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PC EXS</lparam></gate>
<gate>
<ID>794</ID>
<type>DA_FROM</type>
<position>146,-59</position>
<input>
<ID>IN_0</ID>700 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PCDIR</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>72.5,-1</position>
<gparam>LABEL_TEXT Instruction Register and Decode stage 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AM_REGISTER16</type>
<position>33,-50</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>56 </input>
<input>
<ID>IN_10</ID>46 </input>
<input>
<ID>IN_11</ID>44 </input>
<input>
<ID>IN_12</ID>43 </input>
<input>
<ID>IN_13</ID>42 </input>
<input>
<ID>IN_14</ID>41 </input>
<input>
<ID>IN_15</ID>40 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>54 </input>
<input>
<ID>IN_4</ID>52 </input>
<input>
<ID>IN_5</ID>51 </input>
<input>
<ID>IN_6</ID>50 </input>
<input>
<ID>IN_7</ID>49 </input>
<input>
<ID>IN_8</ID>48 </input>
<input>
<ID>IN_9</ID>47 </input>
<output>
<ID>OUT_0</ID>71 </output>
<output>
<ID>OUT_1</ID>72 </output>
<output>
<ID>OUT_10</ID>65 </output>
<output>
<ID>OUT_11</ID>66 </output>
<output>
<ID>OUT_12</ID>59 </output>
<output>
<ID>OUT_13</ID>60 </output>
<output>
<ID>OUT_14</ID>61 </output>
<output>
<ID>OUT_15</ID>58 </output>
<output>
<ID>OUT_2</ID>73 </output>
<output>
<ID>OUT_3</ID>74 </output>
<output>
<ID>OUT_4</ID>67 </output>
<output>
<ID>OUT_5</ID>68 </output>
<output>
<ID>OUT_6</ID>69 </output>
<output>
<ID>OUT_7</ID>70 </output>
<output>
<ID>OUT_8</ID>63 </output>
<output>
<ID>OUT_9</ID>64 </output>
<input>
<ID>clear</ID>37 </input>
<input>
<ID>clock</ID>36 </input>
<input>
<ID>count_enable</ID>38 </input>
<input>
<ID>count_up</ID>38 </input>
<input>
<ID>load</ID>39 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 49156</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>32,-67.5</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>66</ID>
<type>FF_GND</type>
<position>34,-60.5</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>FF_GND</type>
<position>34,-38.5</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>70</ID>
<type>DA_FROM</type>
<position>32,-30.5</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>72</ID>
<type>DA_FROM</type>
<position>9.5,-21</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>73</ID>
<type>DA_FROM</type>
<position>10,-23.5</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>75</ID>
<type>DA_FROM</type>
<position>9.5,-27</position>
<input>
<ID>IN_0</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>76</ID>
<type>DA_FROM</type>
<position>10,-29.5</position>
<input>
<ID>IN_0</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>10,-32.5</position>
<input>
<ID>IN_0</ID>44 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>11,-35</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>79</ID>
<type>DA_FROM</type>
<position>10,-38.5</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>10.5,-41</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>81</ID>
<type>DA_FROM</type>
<position>11.5,-45</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>12,-47.5</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>11,-50.5</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>84</ID>
<type>DA_FROM</type>
<position>12,-53.5</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>664</ID>
<type>AE_DFF_LOW</type>
<position>5,-7.5</position>
<input>
<ID>IN_0</ID>584 </input>
<output>
<ID>OUTINV_0</ID>584 </output>
<output>
<ID>OUT_0</ID>587 </output>
<input>
<ID>clear</ID>583 </input>
<input>
<ID>clock</ID>586 </input>
<input>
<ID>set</ID>585 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>85</ID>
<type>DA_FROM</type>
<position>12,-55.5</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>86</ID>
<type>DA_FROM</type>
<position>12,-58.5</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>666</ID>
<type>EE_VDD</type>
<position>5,-2</position>
<output>
<ID>OUT_0</ID>585 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>87</ID>
<type>DA_FROM</type>
<position>11.5,-61.5</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>88</ID>
<type>DA_FROM</type>
<position>11.5,-65.5</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>668</ID>
<type>EE_VDD</type>
<position>5,-13</position>
<output>
<ID>OUT_0</ID>583 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>669</ID>
<type>DA_FROM</type>
<position>-3.5,-8.5</position>
<input>
<ID>IN_0</ID>586 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>90</ID>
<type>BI_DECODER_4x16</type>
<position>57.5,-26.5</position>
<input>
<ID>ENABLE</ID>62 </input>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>60 </input>
<input>
<ID>IN_2</ID>61 </input>
<input>
<ID>IN_3</ID>58 </input>
<output>
<ID>OUT_12</ID>579 </output>
<output>
<ID>OUT_13</ID>368 </output>
<output>
<ID>OUT_14</ID>261 </output>
<output>
<ID>OUT_15</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>671</ID>
<type>DE_TO</type>
<position>15.5,-8.5</position>
<input>
<ID>IN_0</ID>584 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Execute</lparam></gate>
<gate>
<ID>92</ID>
<type>DA_FROM</type>
<position>46.5,-19</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Execute</lparam></gate>
<gate>
<ID>93</ID>
<type>DE_TO</type>
<position>73.5,-83</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>673</ID>
<type>DE_TO</type>
<position>16.5,-5.5</position>
<input>
<ID>IN_0</ID>587 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>94</ID>
<type>DE_TO</type>
<position>69.5,-83.5</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>95</ID>
<type>DE_TO</type>
<position>66,-84</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>96</ID>
<type>DE_TO</type>
<position>63,-84</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>97</ID>
<type>DE_TO</type>
<position>59.5,-84</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>483</ID>
<type>DE_TO</type>
<position>91.5,-23.5</position>
<input>
<ID>IN_0</ID>579 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MOVEI</lparam></gate>
<gate>
<ID>98</ID>
<type>DE_TO</type>
<position>56,-84</position>
<input>
<ID>IN_0</ID>110 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>291</ID>
<type>DE_TO</type>
<position>92,-14</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID JMP</lparam></gate>
<gate>
<ID>99</ID>
<type>DE_TO</type>
<position>53,-84.5</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>100</ID>
<type>DE_TO</type>
<position>49.5,-84.5</position>
<input>
<ID>IN_0</ID>107 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>293</ID>
<type>DE_TO</type>
<position>148.5,-24.5</position>
<input>
<ID>IN_0</ID>262 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BZ</lparam></gate>
<gate>
<ID>101</ID>
<type>DE_TO</type>
<position>25,-85</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>102</ID>
<type>DE_TO</type>
<position>28.5,-85</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>103</ID>
<type>DE_TO</type>
<position>31.5,-85</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>104</ID>
<type>DE_TO</type>
<position>34.5,-85</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>105</ID>
<type>DE_TO</type>
<position>37.5,-85</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>106</ID>
<type>DE_TO</type>
<position>40,-85</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>107</ID>
<type>DE_TO</type>
<position>42.5,-84.5</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>46,-84.5</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>110</ID>
<type>BI_DECODER_4x16</type>
<position>136.5,-41.5</position>
<input>
<ID>ENABLE</ID>75 </input>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>65 </input>
<input>
<ID>IN_3</ID>66 </input>
<output>
<ID>OUT_13</ID>265 </output>
<output>
<ID>OUT_14</ID>262 </output>
<output>
<ID>OUT_15</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>112</ID>
<type>BI_DECODER_4x16</type>
<position>144,-46</position>
<input>
<ID>ENABLE</ID>76 </input>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>70 </input>
<output>
<ID>OUT_15</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>114</ID>
<type>BI_DECODER_4x16</type>
<position>158.5,-50</position>
<input>
<ID>ENABLE</ID>77 </input>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>116</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>47,-73.5</position>
<input>
<ID>ENABLE_0</ID>125 </input>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_10</ID>65 </input>
<input>
<ID>IN_11</ID>66 </input>
<input>
<ID>IN_12</ID>111 </input>
<input>
<ID>IN_13</ID>111 </input>
<input>
<ID>IN_14</ID>111 </input>
<input>
<ID>IN_15</ID>111 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<input>
<ID>IN_4</ID>67 </input>
<input>
<ID>IN_5</ID>68 </input>
<input>
<ID>IN_6</ID>69 </input>
<input>
<ID>IN_7</ID>70 </input>
<input>
<ID>IN_8</ID>63 </input>
<input>
<ID>IN_9</ID>64 </input>
<output>
<ID>OUT_0</ID>99 </output>
<output>
<ID>OUT_1</ID>100 </output>
<output>
<ID>OUT_10</ID>110 </output>
<output>
<ID>OUT_11</ID>109 </output>
<output>
<ID>OUT_12</ID>98 </output>
<output>
<ID>OUT_13</ID>97 </output>
<output>
<ID>OUT_14</ID>96 </output>
<output>
<ID>OUT_15</ID>95 </output>
<output>
<ID>OUT_2</ID>101 </output>
<output>
<ID>OUT_3</ID>102 </output>
<output>
<ID>OUT_4</ID>103 </output>
<output>
<ID>OUT_5</ID>104 </output>
<output>
<ID>OUT_6</ID>105 </output>
<output>
<ID>OUT_7</ID>106 </output>
<output>
<ID>OUT_8</ID>107 </output>
<output>
<ID>OUT_9</ID>108 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>120</ID>
<type>BA_TRI_STATE</type>
<position>54.5,-67.5</position>
<input>
<ID>ENABLE_0</ID>94 </input>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>111 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>122</ID>
<type>EE_VDD</type>
<position>57.5,-65.5</position>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>126</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>67.5,-60.5</position>
<input>
<ID>ENABLE_0</ID>124 </input>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<output>
<ID>OUT_0</ID>112 </output>
<output>
<ID>OUT_1</ID>113 </output>
<output>
<ID>OUT_2</ID>114 </output>
<output>
<ID>OUT_3</ID>115 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>128</ID>
<type>DE_TO</type>
<position>65,-67.5</position>
<input>
<ID>IN_0</ID>112 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 0</lparam></gate>
<gate>
<ID>129</ID>
<type>DE_TO</type>
<position>67,-67.5</position>
<input>
<ID>IN_0</ID>113 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 1</lparam></gate>
<gate>
<ID>130</ID>
<type>DE_TO</type>
<position>69,-67.5</position>
<input>
<ID>IN_0</ID>114 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 2</lparam></gate>
<gate>
<ID>131</ID>
<type>DE_TO</type>
<position>71,-67.5</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 3</lparam></gate>
<gate>
<ID>132</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>76.5,-60.5</position>
<input>
<ID>ENABLE_0</ID>124 </input>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>70 </input>
<output>
<ID>OUT_0</ID>116 </output>
<output>
<ID>OUT_1</ID>117 </output>
<output>
<ID>OUT_2</ID>118 </output>
<output>
<ID>OUT_3</ID>119 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>133</ID>
<type>DE_TO</type>
<position>74,-67.5</position>
<input>
<ID>IN_0</ID>116 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 4</lparam></gate>
<gate>
<ID>134</ID>
<type>DE_TO</type>
<position>76,-67.5</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 5</lparam></gate>
<gate>
<ID>135</ID>
<type>DE_TO</type>
<position>78,-67.5</position>
<input>
<ID>IN_0</ID>118 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 6</lparam></gate>
<gate>
<ID>136</ID>
<type>DE_TO</type>
<position>80,-67.5</position>
<input>
<ID>IN_0</ID>119 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 7</lparam></gate>
<gate>
<ID>137</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>86,-60.5</position>
<input>
<ID>ENABLE_0</ID>124 </input>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>65 </input>
<input>
<ID>IN_3</ID>66 </input>
<output>
<ID>OUT_0</ID>120 </output>
<output>
<ID>OUT_1</ID>121 </output>
<output>
<ID>OUT_2</ID>122 </output>
<output>
<ID>OUT_3</ID>123 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>138</ID>
<type>DE_TO</type>
<position>83.5,-67.5</position>
<input>
<ID>IN_0</ID>120 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 8</lparam></gate>
<gate>
<ID>139</ID>
<type>DE_TO</type>
<position>85.5,-67.5</position>
<input>
<ID>IN_0</ID>121 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 9</lparam></gate>
<gate>
<ID>140</ID>
<type>DE_TO</type>
<position>87.5,-67.5</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 10</lparam></gate>
<gate>
<ID>141</ID>
<type>DE_TO</type>
<position>89.5,-67.5</position>
<input>
<ID>IN_0</ID>123 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 11</lparam></gate>
<gate>
<ID>143</ID>
<type>DA_FROM</type>
<position>94,-60.5</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID IR-AD</lparam></gate>
<gate>
<ID>145</ID>
<type>DA_FROM</type>
<position>58.5,-73.5</position>
<input>
<ID>IN_0</ID>125 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Imm</lparam></gate>
<gate>
<ID>146</ID>
<type>DE_TO</type>
<position>109.5,-93.5</position>
<input>
<ID>IN_0</ID>126 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Ck2</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_TOGGLE</type>
<position>122,-93.5</position>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>156</ID>
<type>DE_TO</type>
<position>149,-30</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BNZ</lparam></gate>
<gate>
<ID>378</ID>
<type>DE_TO</type>
<position>91.5,-18</position>
<input>
<ID>IN_0</ID>368 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADDI</lparam></gate>
<gate>
<ID>770</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>105,-61</position>
<input>
<ID>ENABLE_0</ID>693 </input>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<output>
<ID>OUT_0</ID>680 </output>
<output>
<ID>OUT_1</ID>681 </output>
<output>
<ID>OUT_2</ID>682 </output>
<output>
<ID>OUT_3</ID>683 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>771</ID>
<type>DE_TO</type>
<position>102.5,-68</position>
<input>
<ID>IN_0</ID>680 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I0</lparam></gate>
<wire>
<ID>579</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62,-23.5,89.5,-23.5</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>62 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>62,-23.5,62,-22</points>
<intersection>-23.5 1</intersection>
<intersection>-22 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>60.5,-22,62,-22</points>
<connection>
<GID>90</GID>
<name>OUT_12</name></connection>
<intersection>62 2</intersection></hsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-12,5,-11.5</points>
<connection>
<GID>664</GID>
<name>clear</name></connection>
<connection>
<GID>668</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>584</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-8.5,11,2.5</points>
<intersection>-8.5 2</intersection>
<intersection>2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,2.5,11,2.5</points>
<intersection>2 3</intersection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-8.5,13.5,-8.5</points>
<connection>
<GID>664</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>671</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>2,-5.5,2,2.5</points>
<connection>
<GID>664</GID>
<name>IN_0</name></connection>
<intersection>2.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>585</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-3.5,5,-3</points>
<connection>
<GID>666</GID>
<name>OUT_0</name></connection>
<connection>
<GID>664</GID>
<name>set</name></connection></vsegment></shape></wire>
<wire>
<ID>586</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-8.5,2,-8.5</points>
<connection>
<GID>669</GID>
<name>IN_0</name></connection>
<intersection>2 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>2,-8.5,2,-8.5</points>
<connection>
<GID>664</GID>
<name>clock</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>587</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8,-5.5,14.5,-5.5</points>
<connection>
<GID>664</GID>
<name>OUT_0</name></connection>
<connection>
<GID>673</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-65.5,32,-59.5</points>
<connection>
<GID>63</GID>
<name>clock</name></connection>
<connection>
<GID>64</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-59.5,34,-59.5</points>
<connection>
<GID>63</GID>
<name>clear</name></connection>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-40.5,34,-39.5</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>-40.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>33,-40.5,34,-40.5</points>
<connection>
<GID>63</GID>
<name>count_up</name></connection>
<connection>
<GID>63</GID>
<name>count_enable</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-40.5,32,-32.5</points>
<connection>
<GID>63</GID>
<name>load</name></connection>
<connection>
<GID>70</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-21,27.5,-21</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>27.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27.5,-42.5,27.5,-21</points>
<intersection>-42.5 4</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>27.5,-42.5,28,-42.5</points>
<connection>
<GID>63</GID>
<name>IN_15</name></connection>
<intersection>27.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-43.5,26,-23.5</points>
<intersection>-43.5 1</intersection>
<intersection>-23.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-43.5,28,-43.5</points>
<connection>
<GID>63</GID>
<name>IN_14</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>12,-23.5,26,-23.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-44.5,24,-27</points>
<intersection>-44.5 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-44.5,28,-44.5</points>
<connection>
<GID>63</GID>
<name>IN_13</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-27,24,-27</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-45.5,22,-29.5</points>
<intersection>-45.5 1</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-45.5,28,-45.5</points>
<connection>
<GID>63</GID>
<name>IN_12</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-29.5,22,-29.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-46.5,21,-32.5</points>
<intersection>-46.5 1</intersection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-46.5,28,-46.5</points>
<connection>
<GID>63</GID>
<name>IN_11</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-32.5,21,-32.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-47.5,20.5,-35</points>
<intersection>-47.5 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-47.5,28,-47.5</points>
<connection>
<GID>63</GID>
<name>IN_10</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-35,20.5,-35</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-48.5,20,-38.5</points>
<intersection>-48.5 1</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-48.5,28,-48.5</points>
<connection>
<GID>63</GID>
<name>IN_9</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-38.5,20,-38.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-49.5,20,-41</points>
<intersection>-49.5 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-49.5,28,-49.5</points>
<connection>
<GID>63</GID>
<name>IN_8</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-41,20,-41</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-50.5,19.5,-45</points>
<intersection>-50.5 1</intersection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-50.5,28,-50.5</points>
<connection>
<GID>63</GID>
<name>IN_7</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-45,19.5,-45</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-51.5,18.5,-47.5</points>
<intersection>-51.5 1</intersection>
<intersection>-47.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-51.5,28,-51.5</points>
<connection>
<GID>63</GID>
<name>IN_6</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-47.5,18.5,-47.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-52.5,17.5,-50.5</points>
<intersection>-52.5 1</intersection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-52.5,28,-52.5</points>
<connection>
<GID>63</GID>
<name>IN_5</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-50.5,17.5,-50.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-53.5,28,-53.5</points>
<connection>
<GID>63</GID>
<name>IN_4</name></connection>
<connection>
<GID>84</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-55.5,23.5,-55.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>23.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>23.5,-55.5,23.5,-54.5</points>
<intersection>-55.5 1</intersection>
<intersection>-54.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>23.5,-54.5,28,-54.5</points>
<connection>
<GID>63</GID>
<name>IN_3</name></connection>
<intersection>23.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-58.5,25,-55.5</points>
<intersection>-58.5 2</intersection>
<intersection>-55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-55.5,28,-55.5</points>
<connection>
<GID>63</GID>
<name>IN_2</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-58.5,25,-58.5</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-61.5,26,-56.5</points>
<intersection>-61.5 2</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-56.5,28,-56.5</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-61.5,26,-61.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-65.5,27.5,-57.5</points>
<intersection>-65.5 2</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-57.5,28,-57.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-65.5,27.5,-65.5</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-31,54.5,-31</points>
<connection>
<GID>90</GID>
<name>IN_3</name></connection>
<intersection>48 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>48,-42.5,48,-31</points>
<intersection>-42.5 5</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>38,-42.5,48,-42.5</points>
<connection>
<GID>63</GID>
<name>OUT_15</name></connection>
<intersection>48 4</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-34,54.5,-34</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>53.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>53.5,-45.5,53.5,-34</points>
<intersection>-45.5 5</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>38,-45.5,53.5,-45.5</points>
<connection>
<GID>63</GID>
<name>OUT_12</name></connection>
<intersection>53.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-33,54.5,-33</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<intersection>51.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51.5,-44.5,51.5,-33</points>
<intersection>-44.5 5</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>38,-44.5,51.5,-44.5</points>
<connection>
<GID>63</GID>
<name>OUT_13</name></connection>
<intersection>51.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-32,54.5,-32</points>
<connection>
<GID>90</GID>
<name>IN_2</name></connection>
<intersection>50 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>50,-43.5,50,-32</points>
<intersection>-43.5 5</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>38,-43.5,50,-43.5</points>
<connection>
<GID>63</GID>
<name>OUT_14</name></connection>
<intersection>50 4</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-19,54.5,-19</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<connection>
<GID>90</GID>
<name>ENABLE</name></connection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-49,133.5,-49</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>38 21</intersection>
<intersection>47.5 13</intersection>
<intersection>84.5 16</intersection>
<intersection>127.5 20</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>47.5,-71.5,47.5,-49</points>
<connection>
<GID>116</GID>
<name>IN_8</name></connection>
<intersection>-49 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>84.5,-58.5,84.5,-49</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>-49 1</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>127.5,-59,127.5,-49</points>
<connection>
<GID>780</GID>
<name>IN_0</name></connection>
<intersection>-49 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>38,-49.5,38,-49</points>
<connection>
<GID>63</GID>
<name>OUT_8</name></connection>
<intersection>-49 1</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-48,133.5,-48</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>38 28</intersection>
<intersection>48.5 13</intersection>
<intersection>85.5 23</intersection>
<intersection>128.5 27</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>48.5,-71.5,48.5,-48</points>
<connection>
<GID>116</GID>
<name>IN_9</name></connection>
<intersection>-48 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>85.5,-58.5,85.5,-48</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<intersection>-48 1</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>128.5,-59,128.5,-48</points>
<connection>
<GID>780</GID>
<name>IN_1</name></connection>
<intersection>-48 1</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>38,-48.5,38,-48</points>
<connection>
<GID>63</GID>
<name>OUT_9</name></connection>
<intersection>-48 1</intersection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-47,133.5,-47</points>
<connection>
<GID>110</GID>
<name>IN_2</name></connection>
<intersection>38 27</intersection>
<intersection>49.5 13</intersection>
<intersection>86.5 22</intersection>
<intersection>129.5 26</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>49.5,-71.5,49.5,-47</points>
<connection>
<GID>116</GID>
<name>IN_10</name></connection>
<intersection>-47 1</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>86.5,-58.5,86.5,-47</points>
<connection>
<GID>137</GID>
<name>IN_2</name></connection>
<intersection>-47 1</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>129.5,-59,129.5,-47</points>
<connection>
<GID>780</GID>
<name>IN_2</name></connection>
<intersection>-47 1</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>38,-47.5,38,-47</points>
<connection>
<GID>63</GID>
<name>OUT_10</name></connection>
<intersection>-47 1</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-46,133.5,-46</points>
<connection>
<GID>110</GID>
<name>IN_3</name></connection>
<intersection>38 32</intersection>
<intersection>50.5 13</intersection>
<intersection>87.5 27</intersection>
<intersection>130.5 31</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>50.5,-71.5,50.5,-46</points>
<connection>
<GID>116</GID>
<name>IN_11</name></connection>
<intersection>-64.5 15</intersection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>50.5,-64.5,54.5,-64.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>50.5 13</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>87.5,-58.5,87.5,-46</points>
<connection>
<GID>137</GID>
<name>IN_3</name></connection>
<intersection>-46 1</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>130.5,-59,130.5,-46</points>
<connection>
<GID>780</GID>
<name>IN_3</name></connection>
<intersection>-46 1</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>38,-46.5,38,-46</points>
<connection>
<GID>63</GID>
<name>OUT_11</name></connection>
<intersection>-46 1</intersection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-53.5,141,-53.5</points>
<connection>
<GID>63</GID>
<name>OUT_4</name></connection>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>43.5 4</intersection>
<intersection>75 8</intersection>
<intersection>112.5 15</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>43.5,-71.5,43.5,-53.5</points>
<connection>
<GID>116</GID>
<name>IN_4</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>75,-58.5,75,-53.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>112.5,-59,112.5,-53.5</points>
<connection>
<GID>775</GID>
<name>IN_0</name></connection>
<intersection>-53.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-20,77,-20</points>
<connection>
<GID>90</GID>
<name>OUT_14</name></connection>
<intersection>77 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77,-20,77,-14</points>
<intersection>-20 1</intersection>
<intersection>-14 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>77,-14,90,-14</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>77 3</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-52.5,141,-52.5</points>
<connection>
<GID>63</GID>
<name>OUT_5</name></connection>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>44.5 4</intersection>
<intersection>76 8</intersection>
<intersection>113.5 15</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>44.5,-71.5,44.5,-52.5</points>
<connection>
<GID>116</GID>
<name>IN_5</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>76,-58.5,76,-52.5</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>113.5,-59,113.5,-52.5</points>
<connection>
<GID>775</GID>
<name>IN_1</name></connection>
<intersection>-52.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140.5,-35,140.5,-24.5</points>
<intersection>-35 4</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>140.5,-24.5,146.5,-24.5</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>140.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>139.5,-35,140.5,-35</points>
<connection>
<GID>110</GID>
<name>OUT_14</name></connection>
<intersection>140.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-51.5,141,-51.5</points>
<connection>
<GID>63</GID>
<name>OUT_6</name></connection>
<connection>
<GID>112</GID>
<name>IN_2</name></connection>
<intersection>45.5 4</intersection>
<intersection>77 8</intersection>
<intersection>114.5 15</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>45.5,-71.5,45.5,-51.5</points>
<connection>
<GID>116</GID>
<name>IN_6</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>77,-58.5,77,-51.5</points>
<connection>
<GID>132</GID>
<name>IN_2</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>114.5,-59,114.5,-51.5</points>
<connection>
<GID>775</GID>
<name>IN_2</name></connection>
<intersection>-51.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-50.5,141,-50.5</points>
<connection>
<GID>63</GID>
<name>OUT_7</name></connection>
<connection>
<GID>112</GID>
<name>IN_3</name></connection>
<intersection>46.5 4</intersection>
<intersection>78 8</intersection>
<intersection>115.5 15</intersection>
<intersection>140.5 16</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>46.5,-71.5,46.5,-50.5</points>
<connection>
<GID>116</GID>
<name>IN_7</name></connection>
<intersection>-50.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>78,-58.5,78,-50.5</points>
<connection>
<GID>132</GID>
<name>IN_3</name></connection>
<intersection>-50.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>115.5,-59,115.5,-50.5</points>
<connection>
<GID>775</GID>
<name>IN_3</name></connection>
<intersection>-50.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>140.5,-60,140.5,-50.5</points>
<connection>
<GID>792</GID>
<name>IN_0</name></connection>
<intersection>-50.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-57.5,155.5,-57.5</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>39.5 7</intersection>
<intersection>66 8</intersection>
<intersection>103.5 12</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>39.5,-71.5,39.5,-57.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>-57.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>66,-58.5,66,-57.5</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-57.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>103.5,-59,103.5,-57.5</points>
<connection>
<GID>770</GID>
<name>IN_0</name></connection>
<intersection>-57.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-36,141,-30</points>
<intersection>-36 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141,-30,147,-30</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139.5,-36,141,-36</points>
<connection>
<GID>110</GID>
<name>OUT_13</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-56.5,155.5,-56.5</points>
<connection>
<GID>63</GID>
<name>OUT_1</name></connection>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>40.5 7</intersection>
<intersection>67 9</intersection>
<intersection>104.5 13</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>40.5,-71.5,40.5,-56.5</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>67,-58.5,67,-56.5</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>104.5,-59,104.5,-56.5</points>
<connection>
<GID>770</GID>
<name>IN_1</name></connection>
<intersection>-56.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-55.5,155.5,-55.5</points>
<connection>
<GID>63</GID>
<name>OUT_2</name></connection>
<connection>
<GID>114</GID>
<name>IN_2</name></connection>
<intersection>41.5 7</intersection>
<intersection>68 8</intersection>
<intersection>105.5 12</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>41.5,-71.5,41.5,-55.5</points>
<connection>
<GID>116</GID>
<name>IN_2</name></connection>
<intersection>-55.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>68,-58.5,68,-55.5</points>
<connection>
<GID>126</GID>
<name>IN_2</name></connection>
<intersection>-55.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>105.5,-59,105.5,-55.5</points>
<connection>
<GID>770</GID>
<name>IN_2</name></connection>
<intersection>-55.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-54.5,155.5,-54.5</points>
<connection>
<GID>63</GID>
<name>OUT_3</name></connection>
<connection>
<GID>114</GID>
<name>IN_3</name></connection>
<intersection>42.5 7</intersection>
<intersection>69 8</intersection>
<intersection>106.5 12</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>42.5,-71.5,42.5,-54.5</points>
<connection>
<GID>116</GID>
<name>IN_3</name></connection>
<intersection>-54.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>69,-58.5,69,-54.5</points>
<connection>
<GID>126</GID>
<name>IN_3</name></connection>
<intersection>-54.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>106.5,-59,106.5,-54.5</points>
<connection>
<GID>770</GID>
<name>IN_3</name></connection>
<intersection>-54.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-34,73.5,-19</points>
<intersection>-34 5</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>60.5,-19,73.5,-19</points>
<connection>
<GID>90</GID>
<name>OUT_15</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>73.5,-34,133.5,-34</points>
<connection>
<GID>110</GID>
<name>ENABLE</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-38.5,140,-34</points>
<intersection>-38.5 3</intersection>
<intersection>-34 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>140,-38.5,141,-38.5</points>
<connection>
<GID>112</GID>
<name>ENABLE</name></connection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>139.5,-34,140,-34</points>
<connection>
<GID>110</GID>
<name>OUT_15</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150.5,-42.5,150.5,-38.5</points>
<intersection>-42.5 1</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-42.5,155.5,-42.5</points>
<connection>
<GID>114</GID>
<name>ENABLE</name></connection>
<intersection>150.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147,-38.5,150.5,-38.5</points>
<connection>
<GID>112</GID>
<name>OUT_15</name></connection>
<intersection>150.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-67.5,57.5,-66.5</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-67.5,57.5,-67.5</points>
<connection>
<GID>120</GID>
<name>ENABLE_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-81,73.5,-75.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>-75.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-75.5,73.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_15</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-81.5,69.5,-76.5</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>-76.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>53.5,-76.5,53.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_14</name></connection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-76.5,69.5,-76.5</points>
<intersection>53.5 1</intersection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-82,66,-77.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>-77.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>52.5,-77.5,52.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_13</name></connection>
<intersection>-77.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>52.5,-77.5,66,-77.5</points>
<intersection>52.5 1</intersection>
<intersection>66 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-82,63,-78</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>-78 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>51.5,-78,51.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_12</name></connection>
<intersection>-78 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-78,63,-78</points>
<intersection>51.5 1</intersection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>25,-83,25,-76</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-76 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>25,-76,39.5,-76</points>
<intersection>25 1</intersection>
<intersection>39.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>39.5,-76,39.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection>
<intersection>-76 2</intersection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-83,28.5,-77</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>-77 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>40.5,-77,40.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_1</name></connection>
<intersection>-77 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-77,40.5,-77</points>
<intersection>28.5 0</intersection>
<intersection>40.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>680</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-66,102.5,-63</points>
<connection>
<GID>771</GID>
<name>IN_0</name></connection>
<intersection>-63 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>102.5,-63,103.5,-63</points>
<connection>
<GID>770</GID>
<name>OUT_0</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-83,31.5,-78</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>-78 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>41.5,-78,41.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_2</name></connection>
<intersection>-78 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-78,41.5,-78</points>
<intersection>31.5 0</intersection>
<intersection>41.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-83,34.5,-78.5</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>-78.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>42.5,-78.5,42.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_3</name></connection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-78.5,42.5,-78.5</points>
<intersection>34.5 0</intersection>
<intersection>42.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>681</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-66,104.5,-63</points>
<connection>
<GID>770</GID>
<name>OUT_1</name></connection>
<connection>
<GID>772</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-83,37.5,-79</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>-79 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>43.5,-79,43.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_4</name></connection>
<intersection>-79 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-79,43.5,-79</points>
<intersection>37.5 0</intersection>
<intersection>43.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>682</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-66,105.5,-63</points>
<connection>
<GID>770</GID>
<name>OUT_2</name></connection>
<intersection>-66 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>105.5,-66,106.5,-66</points>
<connection>
<GID>773</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-83,40,-79.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>-79.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>44.5,-79.5,44.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_5</name></connection>
<intersection>-79.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>40,-79.5,44.5,-79.5</points>
<intersection>40 0</intersection>
<intersection>44.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>683</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-63.5,106.5,-63</points>
<connection>
<GID>770</GID>
<name>OUT_3</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>108.5,-66,108.5,-63.5</points>
<connection>
<GID>774</GID>
<name>IN_0</name></connection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>106.5,-63.5,108.5,-63.5</points>
<intersection>106.5 0</intersection>
<intersection>108.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-82.5,42.5,-80</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>-80 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>45.5,-80,45.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_6</name></connection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-80,45.5,-80</points>
<intersection>42.5 0</intersection>
<intersection>45.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>684</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-66,111.5,-63</points>
<connection>
<GID>776</GID>
<name>IN_0</name></connection>
<intersection>-63 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>111.5,-63,112.5,-63</points>
<connection>
<GID>775</GID>
<name>OUT_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-82.5,46,-79</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-79 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>46.5,-79,46.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_7</name></connection>
<intersection>-79 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>46,-79,46.5,-79</points>
<intersection>46 0</intersection>
<intersection>46.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>685</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-66,113.5,-63</points>
<connection>
<GID>777</GID>
<name>IN_0</name></connection>
<connection>
<GID>775</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-82.5,49.5,-81</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>-81 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>47.5,-81,47.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_8</name></connection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47.5,-81,49.5,-81</points>
<intersection>47.5 1</intersection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>686</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-66,115.5,-64.5</points>
<connection>
<GID>778</GID>
<name>IN_0</name></connection>
<intersection>-64.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>114.5,-64.5,115.5,-64.5</points>
<intersection>114.5 5</intersection>
<intersection>115.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>114.5,-64.5,114.5,-63</points>
<connection>
<GID>775</GID>
<name>OUT_2</name></connection>
<intersection>-64.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-82.5,53,-80</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>-80 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>48.5,-80,48.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_9</name></connection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-80,53,-80</points>
<intersection>48.5 1</intersection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>687</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>117.5,-66,117.5,-63</points>
<connection>
<GID>779</GID>
<name>IN_0</name></connection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>115.5,-63,117.5,-63</points>
<connection>
<GID>775</GID>
<name>OUT_3</name></connection>
<intersection>117.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-82,59.5,-78.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>-78.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>50.5,-78.5,50.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_11</name></connection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-78.5,59.5,-78.5</points>
<intersection>50.5 1</intersection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>688</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-71,124,-65</points>
<connection>
<GID>781</GID>
<name>IN_0</name></connection>
<intersection>-65 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>124,-65,127.5,-65</points>
<intersection>124 0</intersection>
<intersection>127.5 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>127.5,-65,127.5,-63</points>
<connection>
<GID>780</GID>
<name>OUT_0</name></connection>
<intersection>-65 13</intersection></vsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-82,56,-79</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>-79 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>49.5,-79,49.5,-75.5</points>
<connection>
<GID>116</GID>
<name>OUT_10</name></connection>
<intersection>-79 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-79,56,-79</points>
<intersection>49.5 1</intersection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>689</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-66,128.5,-63</points>
<connection>
<GID>780</GID>
<name>OUT_1</name></connection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-66,128.5,-66</points>
<intersection>127 2</intersection>
<intersection>128.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>127,-71,127,-66</points>
<connection>
<GID>782</GID>
<name>IN_0</name></connection>
<intersection>-66 1</intersection></vsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-71.5,54.5,-70</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<connection>
<GID>116</GID>
<name>IN_15</name></connection>
<intersection>-71.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>51.5,-71.5,54.5,-71.5</points>
<connection>
<GID>116</GID>
<name>IN_14</name></connection>
<connection>
<GID>116</GID>
<name>IN_13</name></connection>
<connection>
<GID>116</GID>
<name>IN_12</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>690</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-70.5,129.5,-63</points>
<connection>
<GID>783</GID>
<name>IN_0</name></connection>
<connection>
<GID>780</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-65.5,65,-62.5</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-62.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>65,-62.5,66,-62.5</points>
<connection>
<GID>126</GID>
<name>OUT_0</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-64.5,130.5,-63</points>
<connection>
<GID>780</GID>
<name>OUT_3</name></connection>
<intersection>-64.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>132.5,-71.5,132.5,-64.5</points>
<intersection>-71.5 3</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>130.5,-64.5,132.5,-64.5</points>
<intersection>130.5 0</intersection>
<intersection>132.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>132,-71.5,132.5,-71.5</points>
<connection>
<GID>784</GID>
<name>IN_0</name></connection>
<intersection>132.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-65.5,67,-62.5</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<connection>
<GID>126</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-65.5,69,-62.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-62.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>68,-62.5,69,-62.5</points>
<connection>
<GID>126</GID>
<name>OUT_2</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>693</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-61,117,-61</points>
<connection>
<GID>770</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>775</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>785</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-63,69,-62.5</points>
<connection>
<GID>126</GID>
<name>OUT_3</name></connection>
<intersection>-63 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>71,-65.5,71,-63</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>69,-63,71,-63</points>
<intersection>69 0</intersection>
<intersection>71 1</intersection></hsegment></shape></wire>
<wire>
<ID>694</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-80,136,-72</points>
<connection>
<GID>787</GID>
<name>IN_0</name></connection>
<intersection>-72 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>136,-72,138,-72</points>
<connection>
<GID>786</GID>
<name>OUT_0</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-65.5,74,-62.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>-62.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>74,-62.5,75,-62.5</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>695</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-79.5,139,-72</points>
<connection>
<GID>786</GID>
<name>OUT_1</name></connection>
<connection>
<GID>788</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-65.5,76,-62.5</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<connection>
<GID>132</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>696</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-75,140,-72</points>
<connection>
<GID>786</GID>
<name>OUT_2</name></connection>
<intersection>-75 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>140,-75,143.5,-75</points>
<intersection>140 0</intersection>
<intersection>143.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>143.5,-79,143.5,-75</points>
<connection>
<GID>789</GID>
<name>IN_0</name></connection>
<intersection>-75 6</intersection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-65.5,78,-64</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>-64 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-64,78,-64</points>
<intersection>77 5</intersection>
<intersection>78 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>77,-64,77,-62.5</points>
<connection>
<GID>132</GID>
<name>OUT_2</name></connection>
<intersection>-64 3</intersection></vsegment></shape></wire>
<wire>
<ID>697</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-72.5,141,-72</points>
<connection>
<GID>786</GID>
<name>OUT_3</name></connection>
<intersection>-72.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>147,-79.5,147,-72.5</points>
<connection>
<GID>790</GID>
<name>IN_0</name></connection>
<intersection>-72.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>141,-72.5,147,-72.5</points>
<intersection>141 0</intersection>
<intersection>147 1</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>80,-65.5,80,-62.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>78,-62.5,80,-62.5</points>
<connection>
<GID>132</GID>
<name>OUT_3</name></connection>
<intersection>80 1</intersection></hsegment></shape></wire>
<wire>
<ID>698</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140.5,-66,140.5,-65.5</points>
<connection>
<GID>792</GID>
<name>OUT_0</name></connection>
<intersection>-66 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>138,-66,141,-66</points>
<intersection>138 5</intersection>
<intersection>139 6</intersection>
<intersection>140 7</intersection>
<intersection>140.5 0</intersection>
<intersection>141 8</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>138,-68,138,-66</points>
<connection>
<GID>786</GID>
<name>IN_0</name></connection>
<intersection>-66 4</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>139,-68,139,-66</points>
<connection>
<GID>786</GID>
<name>IN_1</name></connection>
<intersection>-66 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>140,-68,140,-66</points>
<connection>
<GID>786</GID>
<name>IN_2</name></connection>
<intersection>-66 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>141,-68,141,-66</points>
<connection>
<GID>786</GID>
<name>IN_3</name></connection>
<intersection>-66 4</intersection></vsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-65.5,83.5,-62.5</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-62.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>83.5,-62.5,84.5,-62.5</points>
<connection>
<GID>137</GID>
<name>OUT_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>699</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142.5,-70,148,-70</points>
<connection>
<GID>786</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>793</GID>
<name>IN_0</name></connection>
<intersection>143.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>143.5,-70,143.5,-63</points>
<intersection>-70 1</intersection>
<intersection>-63 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>142.5,-63,143.5,-63</points>
<connection>
<GID>792</GID>
<name>ENABLE_0</name></connection>
<intersection>143.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-65.5,85.5,-62.5</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<connection>
<GID>137</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>700</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-61,130,-58.5</points>
<intersection>-61 1</intersection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-61,132,-61</points>
<connection>
<GID>780</GID>
<name>ENABLE_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>130,-58.5,144,-58.5</points>
<intersection>130 0</intersection>
<intersection>144 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>144,-59,144,-58.5</points>
<connection>
<GID>794</GID>
<name>IN_0</name></connection>
<intersection>-58.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-65.5,87.5,-62.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>-62.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>86.5,-62.5,87.5,-62.5</points>
<connection>
<GID>137</GID>
<name>OUT_2</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-63,87.5,-62.5</points>
<connection>
<GID>137</GID>
<name>OUT_3</name></connection>
<intersection>-63 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>89.5,-65.5,89.5,-63</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-63,89.5,-63</points>
<intersection>87.5 0</intersection>
<intersection>89.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-60.5,92,-60.5</points>
<connection>
<GID>132</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>126</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>137</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>143</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56,-73.5,56.5,-73.5</points>
<connection>
<GID>116</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>145</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111.5,-93.5,120,-93.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<connection>
<GID>147</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60.5,-21,89.5,-21</points>
<connection>
<GID>90</GID>
<name>OUT_13</name></connection>
<intersection>89.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>89.5,-21,89.5,-18</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>118.961,-93.7939,435.407,-255.576</PageViewport>
<gate>
<ID>1</ID>
<type>DA_FROM</type>
<position>214,-122</position>
<input>
<ID>IN_0</ID>300 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_AND2</type>
<position>161,-56</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>185 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>DA_FROM</type>
<position>152,-54</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BNZ</lparam></gate>
<gate>
<ID>414</ID>
<type>DE_OR8</type>
<position>132,-255.5</position>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_1</ID>452 </input>
<input>
<ID>IN_2</ID>453 </input>
<input>
<ID>IN_3</ID>454 </input>
<input>
<ID>IN_4</ID>504 </input>
<input>
<ID>IN_5</ID>503 </input>
<input>
<ID>IN_6</ID>502 </input>
<input>
<ID>IN_7</ID>501 </input>
<output>
<ID>OUT</ID>525 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>415</ID>
<type>DA_FROM</type>
<position>121,-243</position>
<input>
<ID>IN_0</ID>451 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MOVEI</lparam></gate>
<gate>
<ID>416</ID>
<type>DA_FROM</type>
<position>111.5,-248.5</position>
<input>
<ID>IN_0</ID>452 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>417</ID>
<type>DA_FROM</type>
<position>112.5,-253.5</position>
<input>
<ID>IN_0</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>444</ID>
<type>DA_FROM</type>
<position>112.5,-256</position>
<input>
<ID>IN_0</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>445</ID>
<type>DE_OR8</type>
<position>132,-221</position>
<input>
<ID>IN_0</ID>526 </input>
<input>
<ID>IN_1</ID>527 </input>
<input>
<ID>IN_2</ID>528 </input>
<input>
<ID>IN_3</ID>529 </input>
<input>
<ID>IN_4</ID>576 </input>
<input>
<ID>IN_5</ID>575 </input>
<input>
<ID>IN_6</ID>574 </input>
<input>
<ID>IN_7</ID>530 </input>
<output>
<ID>OUT</ID>577 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>446</ID>
<type>DA_FROM</type>
<position>112.5,-259</position>
<input>
<ID>IN_0</ID>501 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>447</ID>
<type>DA_FROM</type>
<position>122,-214</position>
<input>
<ID>IN_0</ID>526 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADDI</lparam></gate>
<gate>
<ID>448</ID>
<type>DA_FROM</type>
<position>112.5,-261.5</position>
<input>
<ID>IN_0</ID>502 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>449</ID>
<type>DA_FROM</type>
<position>114,-216.5</position>
<input>
<ID>IN_0</ID>527 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>456</ID>
<type>DA_FROM</type>
<position>113,-264.5</position>
<input>
<ID>IN_0</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>457</ID>
<type>DA_FROM</type>
<position>112.5,-219</position>
<input>
<ID>IN_0</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>458</ID>
<type>DA_FROM</type>
<position>113,-267</position>
<input>
<ID>IN_0</ID>504 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>459</ID>
<type>DA_FROM</type>
<position>112.5,-221.5</position>
<input>
<ID>IN_0</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>460</ID>
<type>DE_TO</type>
<position>144.5,-255.5</position>
<input>
<ID>IN_0</ID>525 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus-Acc</lparam></gate>
<gate>
<ID>461</ID>
<type>DA_FROM</type>
<position>112.5,-224.5</position>
<input>
<ID>IN_0</ID>530 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>463</ID>
<type>DA_FROM</type>
<position>112.5,-227</position>
<input>
<ID>IN_0</ID>574 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>466</ID>
<type>DA_FROM</type>
<position>113,-230</position>
<input>
<ID>IN_0</ID>575 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>468</ID>
<type>DA_FROM</type>
<position>113,-232.5</position>
<input>
<ID>IN_0</ID>576 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>470</ID>
<type>DE_TO</type>
<position>141.5,-221</position>
<input>
<ID>IN_0</ID>577 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Res-Acc</lparam></gate>
<gate>
<ID>113</ID>
<type>DA_FROM</type>
<position>150,-57</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Zero</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>12,-44.5</position>
<gparam>LABEL_TEXT Register Load</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>DE_OR8</type>
<position>33.5,-99.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>195 </input>
<input>
<ID>IN_2</ID>196 </input>
<input>
<ID>IN_3</ID>197 </input>
<input>
<ID>IN_4</ID>201 </input>
<input>
<ID>IN_5</ID>200 </input>
<input>
<ID>IN_6</ID>199 </input>
<input>
<ID>IN_7</ID>198 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>119</ID>
<type>DA_FROM</type>
<position>23.5,-92.5</position>
<input>
<ID>IN_0</ID>194 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADDI</lparam></gate>
<gate>
<ID>121</ID>
<type>DA_FROM</type>
<position>10,-94</position>
<input>
<ID>IN_0</ID>195 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MOVEI</lparam></gate>
<gate>
<ID>123</ID>
<type>DA_FROM</type>
<position>8.5,-97</position>
<input>
<ID>IN_0</ID>196 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>124</ID>
<type>DA_FROM</type>
<position>7.5,-100.5</position>
<input>
<ID>IN_0</ID>197 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>7.5,-103</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>127</ID>
<type>DA_FROM</type>
<position>7.5,-106.5</position>
<input>
<ID>IN_0</ID>199 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>142</ID>
<type>DA_FROM</type>
<position>8,-109.5</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>144</ID>
<type>DA_FROM</type>
<position>8,-114</position>
<input>
<ID>IN_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>149</ID>
<type>DE_TO</type>
<position>43,-99.5</position>
<input>
<ID>IN_0</ID>202 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD Acc</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_LABEL</type>
<position>52,-6</position>
<gparam>LABEL_TEXT Decode stage 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>DE_OR8</type>
<position>133.5,-63.5</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>131 </input>
<input>
<ID>IN_2</ID>133 </input>
<input>
<ID>IN_3</ID>134 </input>
<input>
<ID>IN_4</ID>138 </input>
<input>
<ID>IN_5</ID>137 </input>
<input>
<ID>IN_6</ID>136 </input>
<input>
<ID>IN_7</ID>135 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>153</ID>
<type>AE_SMALL_INVERTER</type>
<position>154.5,-57</position>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>154</ID>
<type>DA_FROM</type>
<position>108,-51</position>
<input>
<ID>IN_0</ID>129 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>157</ID>
<type>DA_FROM</type>
<position>110.5,-55.5</position>
<input>
<ID>IN_0</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>159</ID>
<type>DE_TO</type>
<position>34,-3</position>
<input>
<ID>IN_0</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>161</ID>
<type>FF_GND</type>
<position>30.5,-3</position>
<output>
<ID>OUT_0</ID>132 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>162</ID>
<type>DA_FROM</type>
<position>110,-59.5</position>
<input>
<ID>IN_0</ID>133 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>163</ID>
<type>DA_FROM</type>
<position>110,-63.5</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>164</ID>
<type>DA_FROM</type>
<position>109.5,-66.5</position>
<input>
<ID>IN_0</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_FROM</type>
<position>110.5,-70</position>
<input>
<ID>IN_0</ID>136 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>166</ID>
<type>DA_FROM</type>
<position>111.5,-73.5</position>
<input>
<ID>IN_0</ID>137 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>167</ID>
<type>DA_FROM</type>
<position>111.5,-77.5</position>
<input>
<ID>IN_0</ID>138 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>168</ID>
<type>DE_OR8</type>
<position>325,-65</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>204 </input>
<input>
<ID>IN_2</ID>205 </input>
<input>
<ID>IN_3</ID>206 </input>
<input>
<ID>IN_4</ID>210 </input>
<input>
<ID>IN_5</ID>209 </input>
<input>
<ID>IN_6</ID>208 </input>
<input>
<ID>IN_7</ID>207 </input>
<output>
<ID>OUT</ID>211 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>169</ID>
<type>DE_TO</type>
<position>143,-63.5</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-AD</lparam></gate>
<gate>
<ID>170</ID>
<type>DE_OR8</type>
<position>134.5,-91.5</position>
<input>
<ID>IN_0</ID>140 </input>
<input>
<ID>IN_1</ID>141 </input>
<input>
<ID>IN_2</ID>142 </input>
<input>
<ID>IN_3</ID>143 </input>
<input>
<ID>IN_4</ID>147 </input>
<input>
<ID>IN_5</ID>146 </input>
<input>
<ID>IN_6</ID>145 </input>
<input>
<ID>IN_7</ID>144 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>171</ID>
<type>DA_FROM</type>
<position>121,-82</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADDI</lparam></gate>
<gate>
<ID>172</ID>
<type>DA_FROM</type>
<position>113.5,-85</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MOVEI</lparam></gate>
<gate>
<ID>173</ID>
<type>DA_FROM</type>
<position>111.5,-89.5</position>
<input>
<ID>IN_0</ID>142 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>174</ID>
<type>DA_FROM</type>
<position>111.5,-92.5</position>
<input>
<ID>IN_0</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>175</ID>
<type>DA_FROM</type>
<position>111.5,-95.5</position>
<input>
<ID>IN_0</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>176</ID>
<type>DA_FROM</type>
<position>111.5,-98.5</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>177</ID>
<type>DA_FROM</type>
<position>111.5,-102</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>178</ID>
<type>DA_FROM</type>
<position>111,-107</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>179</ID>
<type>DE_TO</type>
<position>141.5,-91.5</position>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Imm</lparam></gate>
<gate>
<ID>180</ID>
<type>DE_OR8</type>
<position>33.5,-136</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>150 </input>
<input>
<ID>IN_2</ID>151 </input>
<input>
<ID>IN_3</ID>152 </input>
<input>
<ID>IN_4</ID>156 </input>
<input>
<ID>IN_5</ID>155 </input>
<input>
<ID>IN_6</ID>154 </input>
<input>
<ID>IN_7</ID>153 </input>
<output>
<ID>OUT</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>181</ID>
<type>DA_FROM</type>
<position>13.5,-122.5</position>
<input>
<ID>IN_0</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>182</ID>
<type>DA_FROM</type>
<position>13,-127</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>183</ID>
<type>DA_FROM</type>
<position>12.5,-131.5</position>
<input>
<ID>IN_0</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>184</ID>
<type>DA_FROM</type>
<position>12.5,-135.5</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>185</ID>
<type>DA_FROM</type>
<position>12,-139</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>186</ID>
<type>DA_FROM</type>
<position>12,-143.5</position>
<input>
<ID>IN_0</ID>154 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>187</ID>
<type>DA_FROM</type>
<position>12,-147.5</position>
<input>
<ID>IN_0</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>188</ID>
<type>DA_FROM</type>
<position>12,-152</position>
<input>
<ID>IN_0</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>189</ID>
<type>DE_TO</type>
<position>43,-136</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Mem Write</lparam></gate>
<gate>
<ID>190</ID>
<type>DE_OR8</type>
<position>134,-129.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>159 </input>
<input>
<ID>IN_2</ID>160 </input>
<input>
<ID>IN_3</ID>161 </input>
<input>
<ID>IN_4</ID>165 </input>
<input>
<ID>IN_5</ID>164 </input>
<input>
<ID>IN_6</ID>163 </input>
<input>
<ID>IN_7</ID>162 </input>
<output>
<ID>OUT</ID>166 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>579</ID>
<type>DE_OR8</type>
<position>173,-90</position>
<input>
<ID>IN_0</ID>705 </input>
<input>
<ID>IN_1</ID>706 </input>
<input>
<ID>IN_2</ID>707 </input>
<input>
<ID>IN_3</ID>708 </input>
<input>
<ID>IN_4</ID>712 </input>
<input>
<ID>IN_5</ID>711 </input>
<input>
<ID>IN_6</ID>710 </input>
<input>
<ID>IN_7</ID>709 </input>
<output>
<ID>OUT</ID>713 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>191</ID>
<type>DA_FROM</type>
<position>120,-117.5</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>580</ID>
<type>DA_FROM</type>
<position>163,-83</position>
<input>
<ID>IN_0</ID>705 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADDI</lparam></gate>
<gate>
<ID>192</ID>
<type>DA_FROM</type>
<position>115,-122.5</position>
<input>
<ID>IN_0</ID>159 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>581</ID>
<type>DA_FROM</type>
<position>156,-85.5</position>
<input>
<ID>IN_0</ID>706 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>582</ID>
<type>DA_FROM</type>
<position>154.5,-88</position>
<input>
<ID>IN_0</ID>707 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>193</ID>
<type>DA_FROM</type>
<position>114,-127</position>
<input>
<ID>IN_0</ID>160 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>583</ID>
<type>DA_FROM</type>
<position>154.5,-90.5</position>
<input>
<ID>IN_0</ID>708 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>194</ID>
<type>DA_FROM</type>
<position>114,-130.5</position>
<input>
<ID>IN_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>584</ID>
<type>DA_FROM</type>
<position>154.5,-93.5</position>
<input>
<ID>IN_0</ID>709 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>195</ID>
<type>DA_FROM</type>
<position>113.5,-133.5</position>
<input>
<ID>IN_0</ID>162 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>585</ID>
<type>DA_FROM</type>
<position>154.5,-96</position>
<input>
<ID>IN_0</ID>710 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>196</ID>
<type>DA_FROM</type>
<position>113,-136.5</position>
<input>
<ID>IN_0</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>197</ID>
<type>DA_FROM</type>
<position>113,-140</position>
<input>
<ID>IN_0</ID>164 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>587</ID>
<type>DA_FROM</type>
<position>155,-99</position>
<input>
<ID>IN_0</ID>711 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>198</ID>
<type>DA_FROM</type>
<position>114,-143.5</position>
<input>
<ID>IN_0</ID>165 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>199</ID>
<type>DE_TO</type>
<position>143.5,-129.5</position>
<input>
<ID>IN_0</ID>166 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Mem Read</lparam></gate>
<gate>
<ID>200</ID>
<type>DA_FROM</type>
<position>310.5,-51.5</position>
<input>
<ID>IN_0</ID>203 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BRA</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_LABEL</type>
<position>119,-37.5</position>
<gparam>LABEL_TEXT Bus and Memory Controls</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>DA_FROM</type>
<position>304,-57.5</position>
<input>
<ID>IN_0</ID>204 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>204</ID>
<type>DA_FROM</type>
<position>303,-62</position>
<input>
<ID>IN_0</ID>205 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>205</ID>
<type>DA_FROM</type>
<position>304,-65.5</position>
<input>
<ID>IN_0</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>595</ID>
<type>DA_FROM</type>
<position>155,-101.5</position>
<input>
<ID>IN_0</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>206</ID>
<type>DA_FROM</type>
<position>301.5,-68</position>
<input>
<ID>IN_0</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>207</ID>
<type>DA_FROM</type>
<position>303,-71</position>
<input>
<ID>IN_0</ID>208 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>208</ID>
<type>DA_FROM</type>
<position>302,-73.5</position>
<input>
<ID>IN_0</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>598</ID>
<type>DE_TO</type>
<position>188,-90</position>
<input>
<ID>IN_0</ID>713 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID StatEn</lparam></gate>
<gate>
<ID>209</ID>
<type>DA_FROM</type>
<position>302,-79</position>
<input>
<ID>IN_0</ID>210 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>210</ID>
<type>DE_TO</type>
<position>340,-65</position>
<input>
<ID>IN_0</ID>211 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC EXS</lparam></gate>
<gate>
<ID>211</ID>
<type>DE_OR8</type>
<position>33.5,-66.5</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>168 </input>
<input>
<ID>IN_2</ID>169 </input>
<input>
<ID>IN_3</ID>170 </input>
<input>
<ID>IN_4</ID>174 </input>
<input>
<ID>IN_5</ID>173 </input>
<input>
<ID>IN_6</ID>172 </input>
<input>
<ID>IN_7</ID>171 </input>
<output>
<ID>OUT</ID>175 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>212</ID>
<type>DA_FROM</type>
<position>23.5,-56</position>
<input>
<ID>IN_0</ID>167 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID JMP</lparam></gate>
<gate>
<ID>213</ID>
<type>DA_FROM</type>
<position>11,-59.5</position>
<input>
<ID>IN_0</ID>168 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BRA</lparam></gate>
<gate>
<ID>214</ID>
<type>DA_FROM</type>
<position>11,-64</position>
<input>
<ID>IN_0</ID>169 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>215</ID>
<type>DA_FROM</type>
<position>11,-67.5</position>
<input>
<ID>IN_0</ID>170 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>216</ID>
<type>DA_FROM</type>
<position>11,-70.5</position>
<input>
<ID>IN_0</ID>171 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>217</ID>
<type>DA_FROM</type>
<position>11,-74</position>
<input>
<ID>IN_0</ID>172 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>218</ID>
<type>DA_FROM</type>
<position>11.5,-77</position>
<input>
<ID>IN_0</ID>173 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>219</ID>
<type>DA_FROM</type>
<position>11,-82</position>
<input>
<ID>IN_0</ID>174 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>220</ID>
<type>DE_TO</type>
<position>45,-66.5</position>
<input>
<ID>IN_0</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load PC</lparam></gate>
<gate>
<ID>610</ID>
<type>DE_OR8</type>
<position>233.5,-129.5</position>
<input>
<ID>IN_0</ID>300 </input>
<input>
<ID>IN_1</ID>539 </input>
<input>
<ID>IN_2</ID>540 </input>
<input>
<ID>IN_3</ID>541 </input>
<input>
<ID>IN_4</ID>545 </input>
<input>
<ID>IN_5</ID>544 </input>
<input>
<ID>IN_6</ID>543 </input>
<input>
<ID>IN_7</ID>542 </input>
<output>
<ID>OUT</ID>546 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>221</ID>
<type>DE_OR8</type>
<position>324.5,-91.5</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>213 </input>
<input>
<ID>IN_2</ID>214 </input>
<input>
<ID>IN_3</ID>215 </input>
<input>
<ID>IN_4</ID>219 </input>
<input>
<ID>IN_5</ID>218 </input>
<input>
<ID>IN_6</ID>217 </input>
<input>
<ID>IN_7</ID>216 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>222</ID>
<type>DA_FROM</type>
<position>314,-83</position>
<input>
<ID>IN_0</ID>212 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BRA</lparam></gate>
<gate>
<ID>612</ID>
<type>DA_FROM</type>
<position>215.5,-125</position>
<input>
<ID>IN_0</ID>539 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>223</ID>
<type>DA_FROM</type>
<position>305.5,-86.5</position>
<input>
<ID>IN_0</ID>213 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID JMP</lparam></gate>
<gate>
<ID>613</ID>
<type>DA_FROM</type>
<position>214,-127.5</position>
<input>
<ID>IN_0</ID>540 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>224</ID>
<type>DA_FROM</type>
<position>298.5,-89</position>
<input>
<ID>IN_0</ID>214 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>614</ID>
<type>DA_FROM</type>
<position>214,-130</position>
<input>
<ID>IN_0</ID>541 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>225</ID>
<type>DA_FROM</type>
<position>298,-92.5</position>
<input>
<ID>IN_0</ID>215 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>615</ID>
<type>DA_FROM</type>
<position>214,-133</position>
<input>
<ID>IN_0</ID>542 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>226</ID>
<type>DA_FROM</type>
<position>301,-95</position>
<input>
<ID>IN_0</ID>216 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>616</ID>
<type>DA_FROM</type>
<position>214,-135.5</position>
<input>
<ID>IN_0</ID>543 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>227</ID>
<type>DA_FROM</type>
<position>302,-98</position>
<input>
<ID>IN_0</ID>217 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>617</ID>
<type>DA_FROM</type>
<position>214.5,-138.5</position>
<input>
<ID>IN_0</ID>544 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>228</ID>
<type>DA_FROM</type>
<position>302,-102.5</position>
<input>
<ID>IN_0</ID>218 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>618</ID>
<type>DA_FROM</type>
<position>214.5,-141</position>
<input>
<ID>IN_0</ID>545 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>229</ID>
<type>DA_FROM</type>
<position>302.5,-107</position>
<input>
<ID>IN_0</ID>219 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>619</ID>
<type>DE_TO</type>
<position>243,-129.5</position>
<input>
<ID>IN_0</ID>546 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BZero</lparam></gate>
<gate>
<ID>230</ID>
<type>DE_TO</type>
<position>337,-91.5</position>
<input>
<ID>IN_0</ID>220 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-PC</lparam></gate>
<gate>
<ID>231</ID>
<type>DE_OR8</type>
<position>326,-123.5</position>
<input>
<ID>IN_0</ID>221 </input>
<input>
<ID>IN_1</ID>222 </input>
<input>
<ID>IN_2</ID>223 </input>
<input>
<ID>IN_3</ID>224 </input>
<input>
<ID>IN_4</ID>228 </input>
<input>
<ID>IN_5</ID>227 </input>
<input>
<ID>IN_6</ID>226 </input>
<input>
<ID>IN_7</ID>225 </input>
<output>
<ID>OUT</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>621</ID>
<type>AA_LABEL</type>
<position>220,-37.5</position>
<gparam>LABEL_TEXT ALU Controls</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>DA_FROM</type>
<position>312.5,-116</position>
<input>
<ID>IN_0</ID>221 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>622</ID>
<type>DE_OR8</type>
<position>231,-63.5</position>
<input>
<ID>IN_0</ID>547 </input>
<input>
<ID>IN_1</ID>548 </input>
<input>
<ID>IN_2</ID>549 </input>
<input>
<ID>IN_3</ID>550 </input>
<input>
<ID>IN_4</ID>554 </input>
<input>
<ID>IN_5</ID>553 </input>
<input>
<ID>IN_6</ID>552 </input>
<input>
<ID>IN_7</ID>551 </input>
<output>
<ID>OUT</ID>555 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>233</ID>
<type>DA_FROM</type>
<position>308,-119</position>
<input>
<ID>IN_0</ID>222 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID JMP</lparam></gate>
<gate>
<ID>623</ID>
<type>DA_FROM</type>
<position>221,-56.5</position>
<input>
<ID>IN_0</ID>547 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>234</ID>
<type>DA_FROM</type>
<position>306.5,-121.5</position>
<input>
<ID>IN_0</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>624</ID>
<type>DA_FROM</type>
<position>213,-59</position>
<input>
<ID>IN_0</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>235</ID>
<type>DA_FROM</type>
<position>306.5,-124</position>
<input>
<ID>IN_0</ID>224 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>625</ID>
<type>DA_FROM</type>
<position>211.5,-61.5</position>
<input>
<ID>IN_0</ID>549 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>236</ID>
<type>DA_FROM</type>
<position>306.5,-127</position>
<input>
<ID>IN_0</ID>225 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>626</ID>
<type>DA_FROM</type>
<position>211.5,-64</position>
<input>
<ID>IN_0</ID>550 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>237</ID>
<type>DA_FROM</type>
<position>306.5,-129.5</position>
<input>
<ID>IN_0</ID>226 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>627</ID>
<type>DA_FROM</type>
<position>211.5,-67</position>
<input>
<ID>IN_0</ID>551 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>238</ID>
<type>DA_FROM</type>
<position>307,-132.5</position>
<input>
<ID>IN_0</ID>227 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>628</ID>
<type>DA_FROM</type>
<position>211.5,-69.5</position>
<input>
<ID>IN_0</ID>552 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>239</ID>
<type>DA_FROM</type>
<position>307,-135</position>
<input>
<ID>IN_0</ID>228 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>629</ID>
<type>DA_FROM</type>
<position>212,-72.5</position>
<input>
<ID>IN_0</ID>553 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>240</ID>
<type>DE_TO</type>
<position>335.5,-123.5</position>
<input>
<ID>IN_0</ID>229 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCDIR</lparam></gate>
<gate>
<ID>630</ID>
<type>DA_FROM</type>
<position>212,-75</position>
<input>
<ID>IN_0</ID>554 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>241</ID>
<type>AA_LABEL</type>
<position>312,-34.5</position>
<gparam>LABEL_TEXT PC Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>631</ID>
<type>DE_TO</type>
<position>240.5,-63.5</position>
<input>
<ID>IN_0</ID>555 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUBA</lparam></gate>
<gate>
<ID>242</ID>
<type>DE_OR8</type>
<position>326,-145.5</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>231 </input>
<input>
<ID>IN_2</ID>232 </input>
<input>
<ID>IN_3</ID>233 </input>
<input>
<ID>IN_4</ID>237 </input>
<input>
<ID>IN_5</ID>236 </input>
<input>
<ID>IN_6</ID>235 </input>
<input>
<ID>IN_7</ID>234 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>243</ID>
<type>DA_FROM</type>
<position>315.5,-139</position>
<input>
<ID>IN_0</ID>230 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BRA</lparam></gate>
<gate>
<ID>633</ID>
<type>DE_OR8</type>
<position>231,-95</position>
<input>
<ID>IN_0</ID>556 </input>
<input>
<ID>IN_1</ID>557 </input>
<input>
<ID>IN_2</ID>558 </input>
<input>
<ID>IN_3</ID>559 </input>
<input>
<ID>IN_4</ID>563 </input>
<input>
<ID>IN_5</ID>562 </input>
<input>
<ID>IN_6</ID>561 </input>
<input>
<ID>IN_7</ID>560 </input>
<output>
<ID>OUT</ID>564 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>244</ID>
<type>DA_FROM</type>
<position>305,-141.5</position>
<input>
<ID>IN_0</ID>231 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>634</ID>
<type>DA_FROM</type>
<position>221,-88</position>
<input>
<ID>IN_0</ID>556 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>245</ID>
<type>DA_FROM</type>
<position>304,-144</position>
<input>
<ID>IN_0</ID>232 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>635</ID>
<type>DA_FROM</type>
<position>213,-90.5</position>
<input>
<ID>IN_0</ID>557 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>246</ID>
<type>DA_FROM</type>
<position>302.5,-148</position>
<input>
<ID>IN_0</ID>233 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>636</ID>
<type>DA_FROM</type>
<position>211.5,-93</position>
<input>
<ID>IN_0</ID>558 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>247</ID>
<type>DA_FROM</type>
<position>302.5,-150.5</position>
<input>
<ID>IN_0</ID>234 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>637</ID>
<type>DA_FROM</type>
<position>211.5,-95.5</position>
<input>
<ID>IN_0</ID>559 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>248</ID>
<type>DA_FROM</type>
<position>303.5,-152.5</position>
<input>
<ID>IN_0</ID>235 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>638</ID>
<type>DA_FROM</type>
<position>211.5,-98.5</position>
<input>
<ID>IN_0</ID>560 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>249</ID>
<type>DA_FROM</type>
<position>302.5,-156</position>
<input>
<ID>IN_0</ID>236 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>639</ID>
<type>DA_FROM</type>
<position>211.5,-101</position>
<input>
<ID>IN_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>250</ID>
<type>DA_FROM</type>
<position>303.5,-159</position>
<input>
<ID>IN_0</ID>237 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>640</ID>
<type>DA_FROM</type>
<position>212,-104</position>
<input>
<ID>IN_0</ID>562 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>251</ID>
<type>DE_TO</type>
<position>338.5,-145.5</position>
<input>
<ID>IN_0</ID>238 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Offset</lparam></gate>
<gate>
<ID>641</ID>
<type>DA_FROM</type>
<position>212,-106.5</position>
<input>
<ID>IN_0</ID>563 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>252</ID>
<type>DE_OR8</type>
<position>131,-191</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>240 </input>
<input>
<ID>IN_2</ID>241 </input>
<input>
<ID>IN_3</ID>242 </input>
<input>
<ID>IN_4</ID>246 </input>
<input>
<ID>IN_5</ID>245 </input>
<input>
<ID>IN_6</ID>244 </input>
<input>
<ID>IN_7</ID>243 </input>
<output>
<ID>OUT</ID>247 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>642</ID>
<type>DE_TO</type>
<position>240.5,-95</position>
<input>
<ID>IN_0</ID>564 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUBB</lparam></gate>
<gate>
<ID>253</ID>
<type>DA_FROM</type>
<position>120.5,-180</position>
<input>
<ID>IN_0</ID>239 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>643</ID>
<type>DE_OR8</type>
<position>131,-156.5</position>
<input>
<ID>IN_0</ID>565 </input>
<input>
<ID>IN_1</ID>566 </input>
<input>
<ID>IN_2</ID>567 </input>
<input>
<ID>IN_3</ID>568 </input>
<input>
<ID>IN_4</ID>572 </input>
<input>
<ID>IN_5</ID>571 </input>
<input>
<ID>IN_6</ID>570 </input>
<input>
<ID>IN_7</ID>569 </input>
<output>
<ID>OUT</ID>573 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>254</ID>
<type>DA_FROM</type>
<position>108.5,-186.5</position>
<input>
<ID>IN_0</ID>240 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>644</ID>
<type>DA_FROM</type>
<position>120.5,-147</position>
<input>
<ID>IN_0</ID>565 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>645</ID>
<type>DA_FROM</type>
<position>113,-152</position>
<input>
<ID>IN_0</ID>566 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>256</ID>
<type>DA_FROM</type>
<position>107.5,-189.5</position>
<input>
<ID>IN_0</ID>241 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>646</ID>
<type>DA_FROM</type>
<position>111.5,-154.5</position>
<input>
<ID>IN_0</ID>567 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>257</ID>
<type>DA_FROM</type>
<position>106.5,-192</position>
<input>
<ID>IN_0</ID>242 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>647</ID>
<type>DA_FROM</type>
<position>111.5,-157</position>
<input>
<ID>IN_0</ID>568 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>258</ID>
<type>DA_FROM</type>
<position>107,-195</position>
<input>
<ID>IN_0</ID>243 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>648</ID>
<type>DA_FROM</type>
<position>111.5,-160</position>
<input>
<ID>IN_0</ID>569 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>259</ID>
<type>DA_FROM</type>
<position>106.5,-198</position>
<input>
<ID>IN_0</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>649</ID>
<type>DA_FROM</type>
<position>111.5,-162.5</position>
<input>
<ID>IN_0</ID>570 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>260</ID>
<type>DA_FROM</type>
<position>106.5,-200</position>
<input>
<ID>IN_0</ID>245 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>650</ID>
<type>DA_FROM</type>
<position>112,-165.5</position>
<input>
<ID>IN_0</ID>571 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>261</ID>
<type>DA_FROM</type>
<position>106,-204</position>
<input>
<ID>IN_0</ID>246 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>651</ID>
<type>DA_FROM</type>
<position>112,-168</position>
<input>
<ID>IN_0</ID>572 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>262</ID>
<type>DE_TO</type>
<position>142.5,-191</position>
<input>
<ID>IN_0</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-BUS</lparam></gate>
<gate>
<ID>652</ID>
<type>DE_TO</type>
<position>145,-157</position>
<input>
<ID>IN_0</ID>573 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Acc-Bus</lparam></gate>
<gate>
<ID>280</ID>
<type>DE_OR8</type>
<position>326,-168</position>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>253 </input>
<input>
<ID>IN_2</ID>254 </input>
<input>
<ID>IN_3</ID>255 </input>
<input>
<ID>IN_4</ID>259 </input>
<input>
<ID>IN_5</ID>258 </input>
<input>
<ID>IN_6</ID>257 </input>
<input>
<ID>IN_7</ID>256 </input>
<output>
<ID>OUT</ID>260 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>281</ID>
<type>DA_FROM</type>
<position>316,-161</position>
<input>
<ID>IN_0</ID>252 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>282</ID>
<type>DA_FROM</type>
<position>308,-163.5</position>
<input>
<ID>IN_0</ID>253 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>283</ID>
<type>DA_FROM</type>
<position>306.5,-166</position>
<input>
<ID>IN_0</ID>254 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>284</ID>
<type>DA_FROM</type>
<position>306.5,-168.5</position>
<input>
<ID>IN_0</ID>255 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>285</ID>
<type>DA_FROM</type>
<position>306.5,-171.5</position>
<input>
<ID>IN_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>286</ID>
<type>DA_FROM</type>
<position>306.5,-174</position>
<input>
<ID>IN_0</ID>257 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>287</ID>
<type>DA_FROM</type>
<position>307,-177</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>288</ID>
<type>DA_FROM</type>
<position>307,-179.5</position>
<input>
<ID>IN_0</ID>259 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>289</ID>
<type>DE_TO</type>
<position>335.5,-168</position>
<input>
<ID>IN_0</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BUS-PC</lparam></gate>
<gate>
<ID>324</ID>
<type>AA_LABEL</type>
<position>171,-37.5</position>
<gparam>LABEL_TEXT Conditionals</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>325</ID>
<type>DE_OR8</type>
<position>180.5,-61.5</position>
<input>
<ID>IN_0</ID>367 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>339 </input>
<input>
<ID>IN_3</ID>340 </input>
<input>
<ID>IN_4</ID>359 </input>
<input>
<ID>IN_5</ID>358 </input>
<input>
<ID>IN_6</ID>342 </input>
<input>
<ID>IN_7</ID>341 </input>
<output>
<ID>OUT</ID>360 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>326</ID>
<type>DA_FROM</type>
<position>160.5,-47.5</position>
<input>
<ID>IN_0</ID>361 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BZ</lparam></gate>
<gate>
<ID>328</ID>
<type>DA_FROM</type>
<position>159,-60</position>
<input>
<ID>IN_0</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>329</ID>
<type>DA_FROM</type>
<position>159.5,-63</position>
<input>
<ID>IN_0</ID>340 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>330</ID>
<type>DA_FROM</type>
<position>159.5,-66</position>
<input>
<ID>IN_0</ID>341 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>331</ID>
<type>DA_FROM</type>
<position>159.5,-68.5</position>
<input>
<ID>IN_0</ID>342 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>332</ID>
<type>DA_FROM</type>
<position>160,-71.5</position>
<input>
<ID>IN_0</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>333</ID>
<type>DA_FROM</type>
<position>160,-74</position>
<input>
<ID>IN_0</ID>359 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>334</ID>
<type>DE_TO</type>
<position>192.5,-61.5</position>
<input>
<ID>IN_0</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BRA</lparam></gate>
<gate>
<ID>726</ID>
<type>DE_OR8</type>
<position>327,-198</position>
<input>
<ID>IN_0</ID>730 </input>
<input>
<ID>IN_1</ID>731 </input>
<input>
<ID>IN_2</ID>732 </input>
<input>
<ID>IN_3</ID>733 </input>
<input>
<ID>IN_4</ID>737 </input>
<input>
<ID>IN_5</ID>736 </input>
<input>
<ID>IN_6</ID>735 </input>
<input>
<ID>IN_7</ID>734 </input>
<output>
<ID>OUT</ID>738 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>728</ID>
<type>DA_FROM</type>
<position>318.5,-188</position>
<input>
<ID>IN_0</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>730</ID>
<type>DA_FROM</type>
<position>305,-190.5</position>
<input>
<ID>IN_0</ID>731 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>731</ID>
<type>DA_FROM</type>
<position>304,-194.5</position>
<input>
<ID>IN_0</ID>732 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>732</ID>
<type>DA_FROM</type>
<position>303,-198</position>
<input>
<ID>IN_0</ID>733 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>733</ID>
<type>DA_FROM</type>
<position>302,-201</position>
<input>
<ID>IN_0</ID>734 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>738</ID>
<type>DA_FROM</type>
<position>301.5,-205</position>
<input>
<ID>IN_0</ID>735 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>742</ID>
<type>DA_FROM</type>
<position>301.5,-209</position>
<input>
<ID>IN_0</ID>736 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>743</ID>
<type>DA_FROM</type>
<position>301,-214.5</position>
<input>
<ID>IN_0</ID>737 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Low</lparam></gate>
<gate>
<ID>744</ID>
<type>DE_TO</type>
<position>339,-198</position>
<input>
<ID>IN_0</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-ADDR</lparam></gate>
<gate>
<ID>361</ID>
<type>DA_FROM</type>
<position>160.5,-51.5</position>
<input>
<ID>IN_0</ID>366 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Zero</lparam></gate>
<gate>
<ID>365</ID>
<type>AA_AND2</type>
<position>168.5,-50</position>
<input>
<ID>IN_0</ID>361 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>367 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-59,170.5,-56</points>
<intersection>-59 1</intersection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170.5,-59,177.5,-59</points>
<connection>
<GID>325</GID>
<name>IN_1</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>164,-56,170.5,-56</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>170.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-55,155,-54</points>
<intersection>-55 1</intersection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155,-55,158,-55</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-54,155,-54</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-243,129,-243</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<intersection>129 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>129,-252,129,-243</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<intersection>-243 1</intersection></vsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-248.5,127.5,-248.5</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<intersection>127.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>127.5,-253,127.5,-248.5</points>
<intersection>-253 8</intersection>
<intersection>-248.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>127.5,-253,129,-253</points>
<connection>
<GID>414</GID>
<name>IN_1</name></connection>
<intersection>127.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-254,126.5,-253.5</points>
<intersection>-254 1</intersection>
<intersection>-253.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126.5,-254,129,-254</points>
<connection>
<GID>414</GID>
<name>IN_2</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-253.5,126.5,-253.5</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-256,116.5,-255</points>
<intersection>-256 2</intersection>
<intersection>-255 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-255,129,-255</points>
<connection>
<GID>414</GID>
<name>IN_3</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-256,116.5,-256</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-259,117.5,-256</points>
<intersection>-259 2</intersection>
<intersection>-256 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-256,129,-256</points>
<connection>
<GID>414</GID>
<name>IN_7</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-259,117.5,-259</points>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-261.5,119,-257</points>
<intersection>-261.5 2</intersection>
<intersection>-257 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-257,129,-257</points>
<connection>
<GID>414</GID>
<name>IN_6</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-261.5,119,-261.5</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-264.5,121,-258</points>
<intersection>-264.5 2</intersection>
<intersection>-258 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-258,129,-258</points>
<connection>
<GID>414</GID>
<name>IN_5</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-264.5,121,-264.5</points>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-267,123,-259</points>
<intersection>-267 2</intersection>
<intersection>-259 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-259,129,-259</points>
<connection>
<GID>414</GID>
<name>IN_4</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-267,123,-267</points>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>152,-57,152.5,-57</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<connection>
<GID>113</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-51,128,-51</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>128 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128,-60,128,-51</points>
<intersection>-60 5</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>128,-60,130.5,-60</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>128 4</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>112.5,-55.5,126.5,-55.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>126.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>126.5,-61,126.5,-55.5</points>
<intersection>-61 8</intersection>
<intersection>-55.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>126.5,-61,130.5,-61</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<intersection>126.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-3,32,-3</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-62,125.5,-59.5</points>
<intersection>-62 1</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125.5,-62,130.5,-62</points>
<connection>
<GID>152</GID>
<name>IN_2</name></connection>
<intersection>125.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>112,-59.5,125.5,-59.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>125.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>112,-63.5,128,-63.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>128 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128,-63.5,128,-63</points>
<intersection>-63.5 1</intersection>
<intersection>-63 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>128,-63,130.5,-63</points>
<connection>
<GID>152</GID>
<name>IN_3</name></connection>
<intersection>128 3</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-66.5,116.5,-64</points>
<intersection>-66.5 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-64,130.5,-64</points>
<connection>
<GID>152</GID>
<name>IN_7</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-66.5,116.5,-66.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>136,-255.5,142.5,-255.5</points>
<connection>
<GID>414</GID>
<name>OUT</name></connection>
<connection>
<GID>460</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-70,118,-65</points>
<intersection>-70 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-65,130.5,-65</points>
<connection>
<GID>152</GID>
<name>IN_6</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>112.5,-70,118,-70</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-214,129,-214</points>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<intersection>129 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>129,-217.5,129,-214</points>
<connection>
<GID>445</GID>
<name>IN_0</name></connection>
<intersection>-214 1</intersection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-73.5,120,-66</points>
<intersection>-73.5 2</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-66,130.5,-66</points>
<connection>
<GID>152</GID>
<name>IN_5</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-73.5,120,-73.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116,-216.5,127.5,-216.5</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>127.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>127.5,-218.5,127.5,-216.5</points>
<intersection>-218.5 8</intersection>
<intersection>-216.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>127.5,-218.5,129,-218.5</points>
<connection>
<GID>445</GID>
<name>IN_1</name></connection>
<intersection>127.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-77.5,122,-67</points>
<intersection>-77.5 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122,-67,130.5,-67</points>
<connection>
<GID>152</GID>
<name>IN_4</name></connection>
<intersection>122 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-77.5,122,-77.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-219.5,126.5,-219</points>
<intersection>-219.5 1</intersection>
<intersection>-219 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126.5,-219.5,129,-219.5</points>
<connection>
<GID>445</GID>
<name>IN_2</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-219,126.5,-219</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137.5,-63.5,141,-63.5</points>
<connection>
<GID>152</GID>
<name>OUT</name></connection>
<connection>
<GID>169</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-221.5,116.5,-220.5</points>
<intersection>-221.5 2</intersection>
<intersection>-220.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-220.5,129,-220.5</points>
<connection>
<GID>445</GID>
<name>IN_3</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-221.5,116.5,-221.5</points>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-82,129,-82</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>129 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>129,-88,129,-82</points>
<intersection>-88 5</intersection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>129,-88,131.5,-88</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>129 4</intersection></hsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-224.5,117.5,-221.5</points>
<intersection>-224.5 2</intersection>
<intersection>-221.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-221.5,129,-221.5</points>
<connection>
<GID>445</GID>
<name>IN_7</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-224.5,117.5,-224.5</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115.5,-85,127.5,-85</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>127.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>127.5,-89,127.5,-85</points>
<intersection>-89 8</intersection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>127.5,-89,131.5,-89</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>127.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-90,126.5,-89.5</points>
<intersection>-90 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126.5,-90,131.5,-90</points>
<connection>
<GID>170</GID>
<name>IN_2</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-89.5,126.5,-89.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-92.5,116.5,-91</points>
<intersection>-92.5 2</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-91,131.5,-91</points>
<connection>
<GID>170</GID>
<name>IN_3</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-92.5,116.5,-92.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-95.5,117.5,-92</points>
<intersection>-95.5 2</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-92,131.5,-92</points>
<connection>
<GID>170</GID>
<name>IN_7</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-95.5,117.5,-95.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-98.5,119,-93</points>
<intersection>-98.5 2</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-93,131.5,-93</points>
<connection>
<GID>170</GID>
<name>IN_6</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-98.5,119,-98.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-102,121,-94</points>
<intersection>-102 2</intersection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-94,131.5,-94</points>
<connection>
<GID>170</GID>
<name>IN_5</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-102,121,-102</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-107,123,-95</points>
<intersection>-107 2</intersection>
<intersection>-95 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-95,131.5,-95</points>
<connection>
<GID>170</GID>
<name>IN_4</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113,-107,123,-107</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>138.5,-91.5,139.5,-91.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<connection>
<GID>170</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15.5,-122.5,30.5,-122.5</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>30.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>30.5,-132.5,30.5,-122.5</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>-122.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217.5,-125,229,-125</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<intersection>229 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>229,-127,229,-125</points>
<intersection>-127 8</intersection>
<intersection>-125 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>229,-127,230.5,-127</points>
<connection>
<GID>610</GID>
<name>IN_1</name></connection>
<intersection>229 7</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-127,29,-127</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>29 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>29,-133.5,29,-127</points>
<intersection>-133.5 8</intersection>
<intersection>-127 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>29,-133.5,30.5,-133.5</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>29 7</intersection></hsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,-128,228,-127.5</points>
<intersection>-128 1</intersection>
<intersection>-127.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>228,-128,230.5,-128</points>
<connection>
<GID>610</GID>
<name>IN_2</name></connection>
<intersection>228 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-127.5,228,-127.5</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<intersection>228 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-134.5,28,-131.5</points>
<intersection>-134.5 1</intersection>
<intersection>-131.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-134.5,30.5,-134.5</points>
<connection>
<GID>180</GID>
<name>IN_2</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-131.5,28,-131.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-130,218,-129</points>
<intersection>-130 2</intersection>
<intersection>-129 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,-129,230.5,-129</points>
<connection>
<GID>610</GID>
<name>IN_3</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-130,218,-130</points>
<connection>
<GID>614</GID>
<name>IN_0</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14.5,-135.5,30.5,-135.5</points>
<connection>
<GID>180</GID>
<name>IN_3</name></connection>
<connection>
<GID>184</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-133,219,-130</points>
<intersection>-133 2</intersection>
<intersection>-130 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-130,230.5,-130</points>
<connection>
<GID>610</GID>
<name>IN_7</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-133,219,-133</points>
<connection>
<GID>615</GID>
<name>IN_0</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-139,19,-136.5</points>
<intersection>-139 2</intersection>
<intersection>-136.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-136.5,30.5,-136.5</points>
<connection>
<GID>180</GID>
<name>IN_7</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-139,19,-139</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220.5,-135.5,220.5,-131</points>
<intersection>-135.5 2</intersection>
<intersection>-131 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>220.5,-131,230.5,-131</points>
<connection>
<GID>610</GID>
<name>IN_6</name></connection>
<intersection>220.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-135.5,220.5,-135.5</points>
<connection>
<GID>616</GID>
<name>IN_0</name></connection>
<intersection>220.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-143.5,20.5,-137.5</points>
<intersection>-143.5 2</intersection>
<intersection>-137.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-137.5,30.5,-137.5</points>
<connection>
<GID>180</GID>
<name>IN_6</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-143.5,20.5,-143.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222.5,-138.5,222.5,-132</points>
<intersection>-138.5 2</intersection>
<intersection>-132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222.5,-132,230.5,-132</points>
<connection>
<GID>610</GID>
<name>IN_5</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216.5,-138.5,222.5,-138.5</points>
<connection>
<GID>617</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-147.5,22.5,-138.5</points>
<intersection>-147.5 2</intersection>
<intersection>-138.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-138.5,30.5,-138.5</points>
<connection>
<GID>180</GID>
<name>IN_5</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-147.5,22.5,-147.5</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224.5,-141,224.5,-133</points>
<intersection>-141 2</intersection>
<intersection>-133 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224.5,-133,230.5,-133</points>
<connection>
<GID>610</GID>
<name>IN_4</name></connection>
<intersection>224.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216.5,-141,224.5,-141</points>
<connection>
<GID>618</GID>
<name>IN_0</name></connection>
<intersection>224.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-152,24.5,-139.5</points>
<intersection>-152 2</intersection>
<intersection>-139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-139.5,30.5,-139.5</points>
<connection>
<GID>180</GID>
<name>IN_4</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-152,24.5,-152</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>237.5,-129.5,241,-129.5</points>
<connection>
<GID>610</GID>
<name>OUT</name></connection>
<connection>
<GID>619</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-136,41,-136</points>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<connection>
<GID>189</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>223,-56.5,228,-56.5</points>
<connection>
<GID>623</GID>
<name>IN_0</name></connection>
<intersection>228 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>228,-60,228,-56.5</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<intersection>-56.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>122,-117.5,131,-117.5</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>131 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>131,-126,131,-117.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>-117.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215,-59,226.5,-59</points>
<connection>
<GID>624</GID>
<name>IN_0</name></connection>
<intersection>226.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>226.5,-61,226.5,-59</points>
<intersection>-61 8</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>226.5,-61,228,-61</points>
<connection>
<GID>622</GID>
<name>IN_1</name></connection>
<intersection>226.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>117,-122.5,129.5,-122.5</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>129.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>129.5,-127,129.5,-122.5</points>
<intersection>-127 8</intersection>
<intersection>-122.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>129.5,-127,131,-127</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>129.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225.5,-62,225.5,-61.5</points>
<intersection>-62 1</intersection>
<intersection>-61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225.5,-62,228,-62</points>
<connection>
<GID>622</GID>
<name>IN_2</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-61.5,225.5,-61.5</points>
<connection>
<GID>625</GID>
<name>IN_0</name></connection>
<intersection>225.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-128,128.5,-127</points>
<intersection>-128 1</intersection>
<intersection>-127 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128.5,-128,131,-128</points>
<connection>
<GID>190</GID>
<name>IN_2</name></connection>
<intersection>128.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-127,128.5,-127</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>128.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215.5,-64,215.5,-63</points>
<intersection>-64 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215.5,-63,228,-63</points>
<connection>
<GID>622</GID>
<name>IN_3</name></connection>
<intersection>215.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-64,215.5,-64</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>215.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-130.5,118.5,-129</points>
<intersection>-130.5 2</intersection>
<intersection>-129 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118.5,-129,131,-129</points>
<connection>
<GID>190</GID>
<name>IN_3</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-130.5,118.5,-130.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216.5,-67,216.5,-64</points>
<intersection>-67 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216.5,-64,228,-64</points>
<connection>
<GID>622</GID>
<name>IN_7</name></connection>
<intersection>216.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-67,216.5,-67</points>
<connection>
<GID>627</GID>
<name>IN_0</name></connection>
<intersection>216.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-133.5,119.5,-130</points>
<intersection>-133.5 2</intersection>
<intersection>-130 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,-130,131,-130</points>
<connection>
<GID>190</GID>
<name>IN_7</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115.5,-133.5,119.5,-133.5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-69.5,218,-65</points>
<intersection>-69.5 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,-65,228,-65</points>
<connection>
<GID>622</GID>
<name>IN_6</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-69.5,218,-69.5</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-136.5,121,-131</points>
<intersection>-136.5 2</intersection>
<intersection>-131 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-131,131,-131</points>
<connection>
<GID>190</GID>
<name>IN_6</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-136.5,121,-136.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220,-72.5,220,-66</points>
<intersection>-72.5 2</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>220,-66,228,-66</points>
<connection>
<GID>622</GID>
<name>IN_5</name></connection>
<intersection>220 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>214,-72.5,220,-72.5</points>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<intersection>220 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-140,123,-132</points>
<intersection>-140 2</intersection>
<intersection>-132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-132,131,-132</points>
<connection>
<GID>190</GID>
<name>IN_5</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-140,123,-140</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-75,222,-67</points>
<intersection>-75 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222,-67,228,-67</points>
<connection>
<GID>622</GID>
<name>IN_4</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>214,-75,222,-75</points>
<connection>
<GID>630</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-143.5,125,-133</points>
<intersection>-143.5 2</intersection>
<intersection>-133 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-133,131,-133</points>
<connection>
<GID>190</GID>
<name>IN_4</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116,-143.5,125,-143.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235,-63.5,238.5,-63.5</points>
<connection>
<GID>622</GID>
<name>OUT</name></connection>
<connection>
<GID>631</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>138,-129.5,141.5,-129.5</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<connection>
<GID>190</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>223,-88,228,-88</points>
<connection>
<GID>634</GID>
<name>IN_0</name></connection>
<intersection>228 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>228,-91.5,228,-88</points>
<connection>
<GID>633</GID>
<name>IN_0</name></connection>
<intersection>-88 1</intersection></vsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-56,30.5,-56</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>30.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>30.5,-63,30.5,-56</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-56 1</intersection></vsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215,-90.5,226.5,-90.5</points>
<connection>
<GID>635</GID>
<name>IN_0</name></connection>
<intersection>226.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>226.5,-92.5,226.5,-90.5</points>
<intersection>-92.5 8</intersection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>226.5,-92.5,228,-92.5</points>
<connection>
<GID>633</GID>
<name>IN_1</name></connection>
<intersection>226.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-59.5,29,-59.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>29 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>29,-64,29,-59.5</points>
<intersection>-64 8</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>29,-64,30.5,-64</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<intersection>29 7</intersection></hsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225.5,-93.5,225.5,-93</points>
<intersection>-93.5 1</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225.5,-93.5,228,-93.5</points>
<connection>
<GID>633</GID>
<name>IN_2</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-93,225.5,-93</points>
<connection>
<GID>636</GID>
<name>IN_0</name></connection>
<intersection>225.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-65,28,-64</points>
<intersection>-65 1</intersection>
<intersection>-64 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-65,30.5,-65</points>
<connection>
<GID>211</GID>
<name>IN_2</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-64,28,-64</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215.5,-95.5,215.5,-94.5</points>
<intersection>-95.5 2</intersection>
<intersection>-94.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215.5,-94.5,228,-94.5</points>
<connection>
<GID>633</GID>
<name>IN_3</name></connection>
<intersection>215.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-95.5,215.5,-95.5</points>
<connection>
<GID>637</GID>
<name>IN_0</name></connection>
<intersection>215.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-67.5,18,-66</points>
<intersection>-67.5 2</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-66,30.5,-66</points>
<connection>
<GID>211</GID>
<name>IN_3</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-67.5,18,-67.5</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216.5,-98.5,216.5,-95.5</points>
<intersection>-98.5 2</intersection>
<intersection>-95.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216.5,-95.5,228,-95.5</points>
<connection>
<GID>633</GID>
<name>IN_7</name></connection>
<intersection>216.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-98.5,216.5,-98.5</points>
<connection>
<GID>638</GID>
<name>IN_0</name></connection>
<intersection>216.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-70.5,19,-67</points>
<intersection>-70.5 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-67,30.5,-67</points>
<connection>
<GID>211</GID>
<name>IN_7</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-70.5,19,-70.5</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-101,218,-96.5</points>
<intersection>-101 2</intersection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,-96.5,228,-96.5</points>
<connection>
<GID>633</GID>
<name>IN_6</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-101,218,-101</points>
<connection>
<GID>639</GID>
<name>IN_0</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-74,20.5,-68</points>
<intersection>-74 2</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-68,30.5,-68</points>
<connection>
<GID>211</GID>
<name>IN_6</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-74,20.5,-74</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220,-104,220,-97.5</points>
<intersection>-104 2</intersection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>220,-97.5,228,-97.5</points>
<connection>
<GID>633</GID>
<name>IN_5</name></connection>
<intersection>220 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>214,-104,220,-104</points>
<connection>
<GID>640</GID>
<name>IN_0</name></connection>
<intersection>220 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-77,22.5,-69</points>
<intersection>-77 2</intersection>
<intersection>-69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-69,30.5,-69</points>
<connection>
<GID>211</GID>
<name>IN_5</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-77,22.5,-77</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-106.5,222,-98.5</points>
<intersection>-106.5 2</intersection>
<intersection>-98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222,-98.5,228,-98.5</points>
<connection>
<GID>633</GID>
<name>IN_4</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>214,-106.5,222,-106.5</points>
<connection>
<GID>641</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-82,24.5,-70</points>
<intersection>-82 2</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-70,30.5,-70</points>
<connection>
<GID>211</GID>
<name>IN_4</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-82,24.5,-82</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235,-95,238.5,-95</points>
<connection>
<GID>633</GID>
<name>OUT</name></connection>
<connection>
<GID>642</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-66.5,43,-66.5</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<connection>
<GID>220</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>122.5,-147,128,-147</points>
<connection>
<GID>644</GID>
<name>IN_0</name></connection>
<intersection>128 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128,-153,128,-147</points>
<connection>
<GID>643</GID>
<name>IN_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115,-152,126.5,-152</points>
<connection>
<GID>645</GID>
<name>IN_0</name></connection>
<intersection>126.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>126.5,-154,126.5,-152</points>
<intersection>-154 8</intersection>
<intersection>-152 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>126.5,-154,128,-154</points>
<connection>
<GID>643</GID>
<name>IN_1</name></connection>
<intersection>126.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-155,125.5,-154.5</points>
<intersection>-155 1</intersection>
<intersection>-154.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125.5,-155,128,-155</points>
<connection>
<GID>643</GID>
<name>IN_2</name></connection>
<intersection>125.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-154.5,125.5,-154.5</points>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<intersection>125.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-157,115.5,-156</points>
<intersection>-157 2</intersection>
<intersection>-156 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-156,128,-156</points>
<connection>
<GID>643</GID>
<name>IN_3</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-157,115.5,-157</points>
<connection>
<GID>647</GID>
<name>IN_0</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>569</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-160,116.5,-157</points>
<intersection>-160 2</intersection>
<intersection>-157 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-157,128,-157</points>
<connection>
<GID>643</GID>
<name>IN_7</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-160,116.5,-160</points>
<connection>
<GID>648</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-162.5,118,-158</points>
<intersection>-162.5 2</intersection>
<intersection>-158 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-158,128,-158</points>
<connection>
<GID>643</GID>
<name>IN_6</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-162.5,118,-162.5</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-165.5,120,-159</points>
<intersection>-165.5 2</intersection>
<intersection>-159 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-159,128,-159</points>
<connection>
<GID>643</GID>
<name>IN_5</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-165.5,120,-165.5</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-168,122,-160</points>
<intersection>-168 2</intersection>
<intersection>-160 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122,-160,128,-160</points>
<connection>
<GID>643</GID>
<name>IN_4</name></connection>
<intersection>122 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-168,122,-168</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>135,-157,143,-157</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<intersection>135 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>135,-157,135,-156.5</points>
<connection>
<GID>643</GID>
<name>OUT</name></connection>
<intersection>-157 1</intersection></vsegment></shape></wire>
<wire>
<ID>574</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-227,119,-222.5</points>
<intersection>-227 2</intersection>
<intersection>-222.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-222.5,129,-222.5</points>
<connection>
<GID>445</GID>
<name>IN_6</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-227,119,-227</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-57,158,-57</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-230,121,-223.5</points>
<intersection>-230 2</intersection>
<intersection>-223.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-223.5,129,-223.5</points>
<connection>
<GID>445</GID>
<name>IN_5</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-230,121,-230</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-232.5,123,-224.5</points>
<intersection>-232.5 2</intersection>
<intersection>-224.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-224.5,129,-224.5</points>
<connection>
<GID>445</GID>
<name>IN_4</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-232.5,123,-232.5</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>577</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>136,-221,139.5,-221</points>
<connection>
<GID>445</GID>
<name>OUT</name></connection>
<connection>
<GID>470</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-92.5,30.5,-92.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>30.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>30.5,-96,30.5,-92.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>-92.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,-94,29,-94</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>29 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>29,-97,29,-94</points>
<intersection>-97 8</intersection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>29,-97,30.5,-97</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>29 7</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-98,28,-97</points>
<intersection>-98 1</intersection>
<intersection>-97 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-98,30.5,-98</points>
<connection>
<GID>118</GID>
<name>IN_2</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10.5,-97,28,-97</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-100.5,18,-99</points>
<intersection>-100.5 2</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-99,30.5,-99</points>
<connection>
<GID>118</GID>
<name>IN_3</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-100.5,18,-100.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-103,19,-100</points>
<intersection>-103 2</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-100,30.5,-100</points>
<connection>
<GID>118</GID>
<name>IN_7</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-103,19,-103</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-106.5,20.5,-101</points>
<intersection>-106.5 2</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-101,30.5,-101</points>
<connection>
<GID>118</GID>
<name>IN_6</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-106.5,20.5,-106.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-109.5,22.5,-102</points>
<intersection>-109.5 2</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-102,30.5,-102</points>
<connection>
<GID>118</GID>
<name>IN_5</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,-109.5,22.5,-109.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-114,24.5,-103</points>
<intersection>-114 2</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-103,30.5,-103</points>
<connection>
<GID>118</GID>
<name>IN_4</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,-114,24.5,-114</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-99.5,41,-99.5</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<connection>
<GID>149</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>312.5,-51.5,322,-51.5</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>322 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>322,-61.5,322,-51.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>306,-57.5,320.5,-57.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>320.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>320.5,-62.5,320.5,-57.5</points>
<intersection>-62.5 8</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>320.5,-62.5,322,-62.5</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>320.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319.5,-63.5,319.5,-62</points>
<intersection>-63.5 1</intersection>
<intersection>-62 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319.5,-63.5,322,-63.5</points>
<connection>
<GID>168</GID>
<name>IN_2</name></connection>
<intersection>319.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>305,-62,319.5,-62</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>319.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309.5,-65.5,309.5,-64.5</points>
<intersection>-65.5 2</intersection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309.5,-64.5,322,-64.5</points>
<connection>
<GID>168</GID>
<name>IN_3</name></connection>
<intersection>309.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>306,-65.5,309.5,-65.5</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>309.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,-68,310.5,-65.5</points>
<intersection>-68 2</intersection>
<intersection>-65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310.5,-65.5,322,-65.5</points>
<connection>
<GID>168</GID>
<name>IN_7</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-68,310.5,-68</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312,-71,312,-66.5</points>
<intersection>-71 2</intersection>
<intersection>-66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312,-66.5,322,-66.5</points>
<connection>
<GID>168</GID>
<name>IN_6</name></connection>
<intersection>312 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>305,-71,312,-71</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<intersection>312 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314,-73.5,314,-67.5</points>
<intersection>-73.5 2</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,-67.5,322,-67.5</points>
<connection>
<GID>168</GID>
<name>IN_5</name></connection>
<intersection>314 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-73.5,314,-73.5</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>314 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316,-79,316,-68.5</points>
<intersection>-79 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>316,-68.5,322,-68.5</points>
<connection>
<GID>168</GID>
<name>IN_4</name></connection>
<intersection>316 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-79,316,-79</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>316 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>329,-65,338,-65</points>
<connection>
<GID>168</GID>
<name>OUT</name></connection>
<connection>
<GID>210</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>316,-83,321.5,-83</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>321.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>321.5,-88,321.5,-83</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>-83 1</intersection></vsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>307.5,-86.5,320,-86.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>320 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>320,-89,320,-86.5</points>
<intersection>-89 8</intersection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>320,-89,321.5,-89</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>320 7</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319,-90,319,-89</points>
<intersection>-90 1</intersection>
<intersection>-89 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319,-90,321.5,-90</points>
<connection>
<GID>221</GID>
<name>IN_2</name></connection>
<intersection>319 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300.5,-89,319,-89</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>319 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-92.5,309,-91</points>
<intersection>-92.5 2</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309,-91,321.5,-91</points>
<connection>
<GID>221</GID>
<name>IN_3</name></connection>
<intersection>309 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300,-92.5,309,-92.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>309 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,-95,310,-92</points>
<intersection>-95 2</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310,-92,321.5,-92</points>
<connection>
<GID>221</GID>
<name>IN_7</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303,-95,310,-95</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,-98,311.5,-93</points>
<intersection>-98 2</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311.5,-93,321.5,-93</points>
<connection>
<GID>221</GID>
<name>IN_6</name></connection>
<intersection>311.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-98,311.5,-98</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>311.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313.5,-102.5,313.5,-94</points>
<intersection>-102.5 2</intersection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313.5,-94,321.5,-94</points>
<connection>
<GID>221</GID>
<name>IN_5</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-102.5,313.5,-102.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>315.5,-107,315.5,-95</points>
<intersection>-107 2</intersection>
<intersection>-95 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>315.5,-95,321.5,-95</points>
<connection>
<GID>221</GID>
<name>IN_4</name></connection>
<intersection>315.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,-107,315.5,-107</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>315.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>328.5,-91.5,335,-91.5</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<connection>
<GID>230</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>314.5,-116,323,-116</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>323 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>323,-120,323,-116</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>-116 1</intersection></vsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>310,-119,321.5,-119</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>321.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>321.5,-121,321.5,-119</points>
<intersection>-121 8</intersection>
<intersection>-119 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>321.5,-121,323,-121</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<intersection>321.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320.5,-122,320.5,-121.5</points>
<intersection>-122 1</intersection>
<intersection>-121.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320.5,-122,323,-122</points>
<connection>
<GID>231</GID>
<name>IN_2</name></connection>
<intersection>320.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-121.5,320.5,-121.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>320.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,-124,310.5,-123</points>
<intersection>-124 2</intersection>
<intersection>-123 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310.5,-123,323,-123</points>
<connection>
<GID>231</GID>
<name>IN_3</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-124,310.5,-124</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,-127,311.5,-124</points>
<intersection>-127 2</intersection>
<intersection>-124 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311.5,-124,323,-124</points>
<connection>
<GID>231</GID>
<name>IN_7</name></connection>
<intersection>311.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-127,311.5,-127</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>311.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313,-129.5,313,-125</points>
<intersection>-129.5 2</intersection>
<intersection>-125 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313,-125,323,-125</points>
<connection>
<GID>231</GID>
<name>IN_6</name></connection>
<intersection>313 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-129.5,313,-129.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>313 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>315,-132.5,315,-126</points>
<intersection>-132.5 2</intersection>
<intersection>-126 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>315,-126,323,-126</points>
<connection>
<GID>231</GID>
<name>IN_5</name></connection>
<intersection>315 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309,-132.5,315,-132.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>315 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317,-135,317,-127</points>
<intersection>-135 2</intersection>
<intersection>-127 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317,-127,323,-127</points>
<connection>
<GID>231</GID>
<name>IN_4</name></connection>
<intersection>317 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309,-135,317,-135</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>317 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>330,-123.5,333.5,-123.5</points>
<connection>
<GID>231</GID>
<name>OUT</name></connection>
<connection>
<GID>240</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>317.5,-139,322.5,-139</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>322.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>322.5,-142,322.5,-139</points>
<intersection>-142 5</intersection>
<intersection>-139 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>322.5,-142,323,-142</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>322.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>307,-141.5,321,-141.5</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>321 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>321,-143,321,-141.5</points>
<intersection>-143 8</intersection>
<intersection>-141.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>321,-143,323,-143</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>321 7</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>306,-144,323,-144</points>
<connection>
<GID>242</GID>
<name>IN_2</name></connection>
<connection>
<GID>245</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,-148,310,-145</points>
<intersection>-148 2</intersection>
<intersection>-145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310,-145,323,-145</points>
<connection>
<GID>242</GID>
<name>IN_3</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,-148,310,-148</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-150.5,311,-146</points>
<intersection>-150.5 2</intersection>
<intersection>-146 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311,-146,323,-146</points>
<connection>
<GID>242</GID>
<name>IN_7</name></connection>
<intersection>311 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,-150.5,311,-150.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>311 0</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312.5,-152.5,312.5,-147</points>
<intersection>-152.5 2</intersection>
<intersection>-147 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312.5,-147,323,-147</points>
<connection>
<GID>242</GID>
<name>IN_6</name></connection>
<intersection>312.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>305.5,-152.5,312.5,-152.5</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>312.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314.5,-156,314.5,-148</points>
<intersection>-156 2</intersection>
<intersection>-148 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314.5,-148,323,-148</points>
<connection>
<GID>242</GID>
<name>IN_5</name></connection>
<intersection>314.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,-156,314.5,-156</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>314.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316.5,-159,316.5,-149</points>
<intersection>-159 2</intersection>
<intersection>-149 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>316.5,-149,323,-149</points>
<connection>
<GID>242</GID>
<name>IN_4</name></connection>
<intersection>316.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>305.5,-159,316.5,-159</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>316.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>330,-145.5,336.5,-145.5</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<connection>
<GID>242</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>122.5,-180,128,-180</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>128 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128,-187.5,128,-180</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>-180 1</intersection></vsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110.5,-186.5,126.5,-186.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>126.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>126.5,-188.5,126.5,-186.5</points>
<intersection>-188.5 8</intersection>
<intersection>-186.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>126.5,-188.5,128,-188.5</points>
<connection>
<GID>252</GID>
<name>IN_1</name></connection>
<intersection>126.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109.5,-189.5,128,-189.5</points>
<connection>
<GID>252</GID>
<name>IN_2</name></connection>
<connection>
<GID>256</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-192,115.5,-190.5</points>
<intersection>-192 2</intersection>
<intersection>-190.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-190.5,128,-190.5</points>
<connection>
<GID>252</GID>
<name>IN_3</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,-192,115.5,-192</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-195,116.5,-191.5</points>
<intersection>-195 2</intersection>
<intersection>-191.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-191.5,128,-191.5</points>
<connection>
<GID>252</GID>
<name>IN_7</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109,-195,116.5,-195</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-198,118,-192.5</points>
<intersection>-198 2</intersection>
<intersection>-192.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-192.5,128,-192.5</points>
<connection>
<GID>252</GID>
<name>IN_6</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,-198,118,-198</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-200,120,-193.5</points>
<intersection>-200 2</intersection>
<intersection>-193.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-193.5,128,-193.5</points>
<connection>
<GID>252</GID>
<name>IN_5</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,-200,120,-200</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-204,122,-194.5</points>
<intersection>-204 2</intersection>
<intersection>-194.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122,-194.5,128,-194.5</points>
<connection>
<GID>252</GID>
<name>IN_4</name></connection>
<intersection>122 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108,-204,122,-204</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>135,-191,140.5,-191</points>
<connection>
<GID>252</GID>
<name>OUT</name></connection>
<connection>
<GID>262</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>318,-161,323,-161</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>323 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>323,-164.5,323,-161</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>-161 1</intersection></vsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>310,-163.5,321.5,-163.5</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>321.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>321.5,-165.5,321.5,-163.5</points>
<intersection>-165.5 8</intersection>
<intersection>-163.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>321.5,-165.5,323,-165.5</points>
<connection>
<GID>280</GID>
<name>IN_1</name></connection>
<intersection>321.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320.5,-166.5,320.5,-166</points>
<intersection>-166.5 1</intersection>
<intersection>-166 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320.5,-166.5,323,-166.5</points>
<connection>
<GID>280</GID>
<name>IN_2</name></connection>
<intersection>320.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-166,320.5,-166</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>320.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,-168.5,310.5,-167.5</points>
<intersection>-168.5 2</intersection>
<intersection>-167.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310.5,-167.5,323,-167.5</points>
<connection>
<GID>280</GID>
<name>IN_3</name></connection>
<intersection>310.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-168.5,310.5,-168.5</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>310.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,-171.5,311.5,-168.5</points>
<intersection>-171.5 2</intersection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311.5,-168.5,323,-168.5</points>
<connection>
<GID>280</GID>
<name>IN_7</name></connection>
<intersection>311.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-171.5,311.5,-171.5</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>311.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313,-174,313,-169.5</points>
<intersection>-174 2</intersection>
<intersection>-169.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313,-169.5,323,-169.5</points>
<connection>
<GID>280</GID>
<name>IN_6</name></connection>
<intersection>313 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308.5,-174,313,-174</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>313 0</intersection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>315,-177,315,-170.5</points>
<intersection>-177 2</intersection>
<intersection>-170.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>315,-170.5,323,-170.5</points>
<connection>
<GID>280</GID>
<name>IN_5</name></connection>
<intersection>315 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309,-177,315,-177</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>315 0</intersection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317,-179.5,317,-171.5</points>
<intersection>-179.5 2</intersection>
<intersection>-171.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317,-171.5,323,-171.5</points>
<connection>
<GID>280</GID>
<name>IN_4</name></connection>
<intersection>317 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309,-179.5,317,-179.5</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>317 0</intersection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>330,-168,333.5,-168</points>
<connection>
<GID>280</GID>
<name>OUT</name></connection>
<connection>
<GID>289</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-126,230.5,-122</points>
<connection>
<GID>610</GID>
<name>IN_0</name></connection>
<intersection>-122 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216,-122,230.5,-122</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>230.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>705</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165,-83,170,-83</points>
<connection>
<GID>580</GID>
<name>IN_0</name></connection>
<intersection>170 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>170,-86.5,170,-83</points>
<connection>
<GID>579</GID>
<name>IN_0</name></connection>
<intersection>-83 1</intersection></vsegment></shape></wire>
<wire>
<ID>706</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>158,-85.5,168.5,-85.5</points>
<connection>
<GID>581</GID>
<name>IN_0</name></connection>
<intersection>168.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>168.5,-87.5,168.5,-85.5</points>
<intersection>-87.5 8</intersection>
<intersection>-85.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>168.5,-87.5,170,-87.5</points>
<connection>
<GID>579</GID>
<name>IN_1</name></connection>
<intersection>168.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>707</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-88.5,167.5,-88</points>
<intersection>-88.5 1</intersection>
<intersection>-88 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167.5,-88.5,170,-88.5</points>
<connection>
<GID>579</GID>
<name>IN_2</name></connection>
<intersection>167.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-88,167.5,-88</points>
<connection>
<GID>582</GID>
<name>IN_0</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>708</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,-90.5,157.5,-89.5</points>
<intersection>-90.5 3</intersection>
<intersection>-89.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-89.5,170,-89.5</points>
<connection>
<GID>579</GID>
<name>IN_3</name></connection>
<intersection>157.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>156.5,-90.5,157.5,-90.5</points>
<connection>
<GID>583</GID>
<name>IN_0</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>709</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158.5,-93.5,158.5,-90.5</points>
<intersection>-93.5 2</intersection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158.5,-90.5,170,-90.5</points>
<connection>
<GID>579</GID>
<name>IN_7</name></connection>
<intersection>158.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-93.5,158.5,-93.5</points>
<connection>
<GID>584</GID>
<name>IN_0</name></connection>
<intersection>158.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>710</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-96,160,-91.5</points>
<intersection>-96 2</intersection>
<intersection>-91.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160,-91.5,170,-91.5</points>
<connection>
<GID>579</GID>
<name>IN_6</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-96,160,-96</points>
<connection>
<GID>585</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment></shape></wire>
<wire>
<ID>711</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-99,162,-92.5</points>
<intersection>-99 2</intersection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162,-92.5,170,-92.5</points>
<connection>
<GID>579</GID>
<name>IN_5</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157,-99,162,-99</points>
<connection>
<GID>587</GID>
<name>IN_0</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>712</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164,-101.5,164,-93.5</points>
<intersection>-101.5 2</intersection>
<intersection>-93.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>164,-93.5,170,-93.5</points>
<connection>
<GID>579</GID>
<name>IN_4</name></connection>
<intersection>164 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157,-101.5,164,-101.5</points>
<connection>
<GID>595</GID>
<name>IN_0</name></connection>
<intersection>164 0</intersection></hsegment></shape></wire>
<wire>
<ID>713</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-90,186,-90</points>
<connection>
<GID>579</GID>
<name>OUT</name></connection>
<connection>
<GID>598</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161,-60,177.5,-60</points>
<connection>
<GID>325</GID>
<name>IN_2</name></connection>
<connection>
<GID>328</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-63,165,-61</points>
<intersection>-63 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165,-61,177.5,-61</points>
<connection>
<GID>325</GID>
<name>IN_3</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161.5,-63,165,-63</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>730</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>320.5,-188,324,-188</points>
<connection>
<GID>728</GID>
<name>IN_0</name></connection>
<intersection>324 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>324,-194.5,324,-188</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<intersection>-188 1</intersection></vsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-66,166,-62</points>
<intersection>-66 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-62,177.5,-62</points>
<connection>
<GID>325</GID>
<name>IN_7</name></connection>
<intersection>166 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161.5,-66,166,-66</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>731</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>307,-190.5,322.5,-190.5</points>
<connection>
<GID>730</GID>
<name>IN_0</name></connection>
<intersection>322.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>322.5,-195.5,322.5,-190.5</points>
<intersection>-195.5 8</intersection>
<intersection>-190.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>322.5,-195.5,324,-195.5</points>
<connection>
<GID>726</GID>
<name>IN_1</name></connection>
<intersection>322.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-68.5,167.5,-63</points>
<intersection>-68.5 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167.5,-63,177.5,-63</points>
<connection>
<GID>325</GID>
<name>IN_6</name></connection>
<intersection>167.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161.5,-68.5,167.5,-68.5</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>732</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321.5,-196.5,321.5,-194.5</points>
<intersection>-196.5 1</intersection>
<intersection>-194.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321.5,-196.5,324,-196.5</points>
<connection>
<GID>726</GID>
<name>IN_2</name></connection>
<intersection>321.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>306,-194.5,321.5,-194.5</points>
<connection>
<GID>731</GID>
<name>IN_0</name></connection>
<intersection>321.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>733</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>305,-198,324,-198</points>
<connection>
<GID>732</GID>
<name>IN_0</name></connection>
<intersection>324 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>324,-198,324,-197.5</points>
<connection>
<GID>726</GID>
<name>IN_3</name></connection>
<intersection>-198 1</intersection></vsegment></shape></wire>
<wire>
<ID>734</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312.5,-201,312.5,-198.5</points>
<intersection>-201 2</intersection>
<intersection>-198.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312.5,-198.5,324,-198.5</points>
<connection>
<GID>726</GID>
<name>IN_7</name></connection>
<intersection>312.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-201,312.5,-201</points>
<connection>
<GID>733</GID>
<name>IN_0</name></connection>
<intersection>312.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>735</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314,-205,314,-199.5</points>
<intersection>-205 2</intersection>
<intersection>-199.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,-199.5,324,-199.5</points>
<connection>
<GID>726</GID>
<name>IN_6</name></connection>
<intersection>314 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-205,314,-205</points>
<connection>
<GID>738</GID>
<name>IN_0</name></connection>
<intersection>314 0</intersection></hsegment></shape></wire>
<wire>
<ID>736</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316,-209,316,-200.5</points>
<intersection>-209 2</intersection>
<intersection>-200.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>316,-200.5,324,-200.5</points>
<connection>
<GID>726</GID>
<name>IN_5</name></connection>
<intersection>316 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-209,316,-209</points>
<connection>
<GID>742</GID>
<name>IN_0</name></connection>
<intersection>316 0</intersection></hsegment></shape></wire>
<wire>
<ID>737</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>318,-214.5,318,-201.5</points>
<intersection>-214.5 2</intersection>
<intersection>-201.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318,-201.5,324,-201.5</points>
<connection>
<GID>726</GID>
<name>IN_4</name></connection>
<intersection>318 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303,-214.5,318,-214.5</points>
<connection>
<GID>743</GID>
<name>IN_0</name></connection>
<intersection>318 0</intersection></hsegment></shape></wire>
<wire>
<ID>738</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>331,-198,337,-198</points>
<connection>
<GID>726</GID>
<name>OUT</name></connection>
<connection>
<GID>744</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-71.5,169.5,-64</points>
<intersection>-71.5 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-64,177.5,-64</points>
<connection>
<GID>325</GID>
<name>IN_5</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162,-71.5,169.5,-71.5</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171.5,-74,171.5,-65</points>
<intersection>-74 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171.5,-65,177.5,-65</points>
<connection>
<GID>325</GID>
<name>IN_4</name></connection>
<intersection>171.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162,-74,171.5,-74</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>171.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>184.5,-61.5,190.5,-61.5</points>
<connection>
<GID>325</GID>
<name>OUT</name></connection>
<connection>
<GID>334</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-49,163.5,-47.5</points>
<intersection>-49 1</intersection>
<intersection>-47.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163.5,-49,165.5,-49</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-47.5,163.5,-47.5</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-51.5,163.5,-51</points>
<intersection>-51.5 2</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163.5,-51,165.5,-51</points>
<connection>
<GID>365</GID>
<name>IN_1</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-51.5,163.5,-51.5</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-58,174,-50</points>
<intersection>-58 1</intersection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174,-58,177.5,-58</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>171.5,-50,174,-50</points>
<connection>
<GID>365</GID>
<name>OUT</name></connection>
<intersection>174 0</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-126.638,140.156,623.456,-243.328</PageViewport>
<gate>
<ID>389</ID>
<type>GA_LED</type>
<position>-113.5,-5.5</position>
<input>
<ID>N_in2</ID>315 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>390</ID>
<type>DE_TO</type>
<position>-122,-97.5</position>
<input>
<ID>IN_0</ID>661 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A12</lparam></gate>
<gate>
<ID>391</ID>
<type>DE_TO</type>
<position>-127.5,-96</position>
<input>
<ID>IN_0</ID>334 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A13</lparam></gate>
<gate>
<ID>392</ID>
<type>DE_TO</type>
<position>-121,-94.5</position>
<input>
<ID>IN_0</ID>335 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A14</lparam></gate>
<gate>
<ID>393</ID>
<type>DE_TO</type>
<position>-127,-93</position>
<input>
<ID>IN_0</ID>336 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A15</lparam></gate>
<gate>
<ID>394</ID>
<type>DE_TO</type>
<position>-117,-8.5</position>
<input>
<ID>IN_0</ID>315 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Zero</lparam></gate>
<gate>
<ID>395</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>-54,-44</position>
<input>
<ID>ENABLE_0</ID>396 </input>
<input>
<ID>IN_0</ID>350 </input>
<input>
<ID>IN_1</ID>349 </input>
<input>
<ID>IN_2</ID>348 </input>
<input>
<ID>IN_3</ID>347 </input>
<output>
<ID>OUT_0</ID>346 </output>
<output>
<ID>OUT_1</ID>345 </output>
<output>
<ID>OUT_2</ID>344 </output>
<output>
<ID>OUT_3</ID>343 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>396</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>-50.5,-34.5</position>
<input>
<ID>ENABLE_0</ID>369 </input>
<input>
<ID>IN_0</ID>354 </input>
<input>
<ID>IN_1</ID>353 </input>
<input>
<ID>IN_2</ID>352 </input>
<input>
<ID>IN_3</ID>351 </input>
<output>
<ID>OUT_0</ID>343 </output>
<output>
<ID>OUT_1</ID>344 </output>
<output>
<ID>OUT_2</ID>345 </output>
<output>
<ID>OUT_3</ID>346 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>397</ID>
<type>BE_NOR4</type>
<position>-88.5,-84.5</position>
<input>
<ID>IN_0</ID>661 </input>
<input>
<ID>IN_1</ID>334 </input>
<input>
<ID>IN_2</ID>335 </input>
<input>
<ID>IN_3</ID>336 </input>
<output>
<ID>OUT</ID>418 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>398</ID>
<type>DA_FROM</type>
<position>-61,-42.5</position>
<input>
<ID>IN_0</ID>347 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A15</lparam></gate>
<gate>
<ID>399</ID>
<type>DA_FROM</type>
<position>-65.5,-43.5</position>
<input>
<ID>IN_0</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A14</lparam></gate>
<gate>
<ID>400</ID>
<type>DA_FROM</type>
<position>-71,-44.5</position>
<input>
<ID>IN_0</ID>349 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A13</lparam></gate>
<gate>
<ID>401</ID>
<type>DA_FROM</type>
<position>-77,-45.5</position>
<input>
<ID>IN_0</ID>350 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A12</lparam></gate>
<gate>
<ID>402</ID>
<type>DA_FROM</type>
<position>-2,-23.5</position>
<input>
<ID>IN_0</ID>351 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>403</ID>
<type>DA_FROM</type>
<position>-6,-23</position>
<input>
<ID>IN_0</ID>352 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>404</ID>
<type>DA_FROM</type>
<position>-10,-22.5</position>
<input>
<ID>IN_0</ID>353 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>405</ID>
<type>DA_FROM</type>
<position>-13,-22.5</position>
<input>
<ID>IN_0</ID>354 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>406</ID>
<type>DA_FROM</type>
<position>-49.5,-50</position>
<input>
<ID>IN_0</ID>355 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>407</ID>
<type>FF_GND</type>
<position>-42,-49.5</position>
<output>
<ID>OUT_0</ID>356 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>408</ID>
<type>FF_GND</type>
<position>-43,-36.5</position>
<output>
<ID>OUT_0</ID>357 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>409</ID>
<type>DA_FROM</type>
<position>101.5,-25</position>
<input>
<ID>IN_0</ID>397 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Res-Acc</lparam></gate>
<gate>
<ID>410</ID>
<type>DA_FROM</type>
<position>244.5,-31.5</position>
<input>
<ID>IN_0</ID>398 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Res-Acc</lparam></gate>
<gate>
<ID>411</ID>
<type>DA_FROM</type>
<position>387,-28.5</position>
<input>
<ID>IN_0</ID>450 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Res-Acc</lparam></gate>
<gate>
<ID>418</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>101.5,-44.5</position>
<input>
<ID>ENABLE_0</ID>397 </input>
<input>
<ID>IN_0</ID>406 </input>
<input>
<ID>IN_1</ID>405 </input>
<input>
<ID>IN_2</ID>404 </input>
<input>
<ID>IN_3</ID>403 </input>
<output>
<ID>OUT_0</ID>402 </output>
<output>
<ID>OUT_1</ID>401 </output>
<output>
<ID>OUT_2</ID>400 </output>
<output>
<ID>OUT_3</ID>399 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>419</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>105,-35</position>
<input>
<ID>ENABLE_0</ID>370 </input>
<input>
<ID>IN_0</ID>410 </input>
<input>
<ID>IN_1</ID>409 </input>
<input>
<ID>IN_2</ID>408 </input>
<input>
<ID>IN_3</ID>407 </input>
<output>
<ID>OUT_0</ID>399 </output>
<output>
<ID>OUT_1</ID>400 </output>
<output>
<ID>OUT_2</ID>401 </output>
<output>
<ID>OUT_3</ID>402 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>420</ID>
<type>DA_FROM</type>
<position>94.5,-43</position>
<input>
<ID>IN_0</ID>403 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A11</lparam></gate>
<gate>
<ID>421</ID>
<type>DA_FROM</type>
<position>90,-44</position>
<input>
<ID>IN_0</ID>404 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A10</lparam></gate>
<gate>
<ID>422</ID>
<type>DA_FROM</type>
<position>84.5,-45</position>
<input>
<ID>IN_0</ID>405 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A9</lparam></gate>
<gate>
<ID>423</ID>
<type>DA_FROM</type>
<position>78.5,-46</position>
<input>
<ID>IN_0</ID>406 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A8</lparam></gate>
<gate>
<ID>424</ID>
<type>DA_FROM</type>
<position>156,-25</position>
<input>
<ID>IN_0</ID>407 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>425</ID>
<type>DA_FROM</type>
<position>152,-24.5</position>
<input>
<ID>IN_0</ID>408 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>426</ID>
<type>DA_FROM</type>
<position>148,-24</position>
<input>
<ID>IN_0</ID>409 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>427</ID>
<type>DA_FROM</type>
<position>145,-24</position>
<input>
<ID>IN_0</ID>410 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>428</ID>
<type>DA_FROM</type>
<position>106,-50.5</position>
<input>
<ID>IN_0</ID>411 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>429</ID>
<type>FF_GND</type>
<position>113.5,-50</position>
<output>
<ID>OUT_0</ID>412 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>430</ID>
<type>FF_GND</type>
<position>112.5,-37.5</position>
<output>
<ID>OUT_0</ID>413 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>431</ID>
<type>AE_FULLADDER_4BIT</type>
<position>118,-89.5</position>
<input>
<ID>IN_0</ID>380 </input>
<input>
<ID>IN_1</ID>382 </input>
<input>
<ID>IN_2</ID>383 </input>
<input>
<ID>IN_3</ID>384 </input>
<input>
<ID>IN_B_0</ID>362 </input>
<input>
<ID>IN_B_1</ID>363 </input>
<input>
<ID>IN_B_2</ID>364 </input>
<input>
<ID>IN_B_3</ID>365 </input>
<output>
<ID>OUT_0</ID>390 </output>
<output>
<ID>OUT_1</ID>391 </output>
<output>
<ID>OUT_2</ID>392 </output>
<output>
<ID>OUT_3</ID>393 </output>
<input>
<ID>carry_in</ID>523 </input>
<output>
<ID>carry_out</ID>414 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>432</ID>
<type>AI_XOR2</type>
<position>139,-68</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>375 </input>
<output>
<ID>OUT</ID>362 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>433</ID>
<type>AI_XOR2</type>
<position>132.5,-68</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>376 </input>
<output>
<ID>OUT</ID>363 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>434</ID>
<type>AI_XOR2</type>
<position>127,-68</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>377 </input>
<output>
<ID>OUT</ID>364 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>435</ID>
<type>AI_XOR2</type>
<position>120,-68</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>378 </input>
<output>
<ID>OUT</ID>365 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>436</ID>
<type>DA_FROM</type>
<position>114,-61</position>
<input>
<ID>IN_0</ID>374 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>437</ID>
<type>DA_FROM</type>
<position>107.5,-60.5</position>
<input>
<ID>IN_0</ID>373 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>438</ID>
<type>DA_FROM</type>
<position>102.5,-60</position>
<input>
<ID>IN_0</ID>372 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>439</ID>
<type>DA_FROM</type>
<position>96,-60</position>
<input>
<ID>IN_0</ID>371 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>440</ID>
<type>AI_XOR2</type>
<position>115,-69</position>
<input>
<ID>IN_0</ID>388 </input>
<input>
<ID>IN_1</ID>374 </input>
<output>
<ID>OUT</ID>379 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>441</ID>
<type>AI_XOR2</type>
<position>108.5,-69</position>
<input>
<ID>IN_0</ID>388 </input>
<input>
<ID>IN_1</ID>373 </input>
<output>
<ID>OUT</ID>381 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>442</ID>
<type>AI_XOR2</type>
<position>103.5,-69</position>
<input>
<ID>IN_0</ID>388 </input>
<input>
<ID>IN_1</ID>372 </input>
<output>
<ID>OUT</ID>385 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>443</ID>
<type>AI_XOR2</type>
<position>97,-69</position>
<input>
<ID>IN_0</ID>388 </input>
<input>
<ID>IN_1</ID>371 </input>
<output>
<ID>OUT</ID>386 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>450</ID>
<type>AA_REGISTER4</type>
<position>112.5,-45</position>
<input>
<ID>IN_0</ID>402 </input>
<input>
<ID>IN_1</ID>401 </input>
<input>
<ID>IN_2</ID>400 </input>
<input>
<ID>IN_3</ID>399 </input>
<output>
<ID>OUT_0</ID>375 </output>
<output>
<ID>OUT_1</ID>376 </output>
<output>
<ID>OUT_2</ID>377 </output>
<output>
<ID>OUT_3</ID>378 </output>
<input>
<ID>clear</ID>412 </input>
<input>
<ID>clock</ID>411 </input>
<input>
<ID>count_enable</ID>413 </input>
<input>
<ID>count_up</ID>413 </input>
<input>
<ID>load</ID>415 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>451</ID>
<type>AA_AND2</type>
<position>116,-77.5</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>380 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>452</ID>
<type>AA_AND2</type>
<position>109.5,-78</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>381 </input>
<output>
<ID>OUT</ID>382 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>453</ID>
<type>AA_AND2</type>
<position>104.5,-78</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>385 </input>
<output>
<ID>OUT</ID>383 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>454</ID>
<type>AA_AND2</type>
<position>98,-78</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>386 </input>
<output>
<ID>OUT</ID>384 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>455</ID>
<type>AE_SMALL_INVERTER</type>
<position>93.5,-73.5</position>
<input>
<ID>IN_0</ID>416 </input>
<output>
<ID>OUT_0</ID>387 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>462</ID>
<type>DA_FROM</type>
<position>122.5,-36</position>
<input>
<ID>IN_0</ID>415 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LD Acc</lparam></gate>
<gate>
<ID>464</ID>
<type>DA_FROM</type>
<position>84.5,-73.5</position>
<input>
<ID>IN_0</ID>416 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BZero</lparam></gate>
<gate>
<ID>465</ID>
<type>DA_FROM</type>
<position>-68.5,-69.5</position>
<input>
<ID>IN_0</ID>417 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BZero</lparam></gate>
<gate>
<ID>467</ID>
<type>DE_TO</type>
<position>-88.5,-62</position>
<input>
<ID>IN_0</ID>418 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z15-12</lparam></gate>
<gate>
<ID>471</ID>
<type>DA_FROM</type>
<position>-116.5,-37</position>
<input>
<ID>IN_0</ID>624 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z15-12</lparam></gate>
<gate>
<ID>472</ID>
<type>DA_FROM</type>
<position>-113.5,-37</position>
<input>
<ID>IN_0</ID>625 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z11-8</lparam></gate>
<gate>
<ID>475</ID>
<type>DE_TO</type>
<position>66.5,-98</position>
<input>
<ID>IN_0</ID>390 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A8</lparam></gate>
<gate>
<ID>476</ID>
<type>DE_TO</type>
<position>61,-96.5</position>
<input>
<ID>IN_0</ID>391 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A9</lparam></gate>
<gate>
<ID>477</ID>
<type>DE_TO</type>
<position>67.5,-95</position>
<input>
<ID>IN_0</ID>392 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A10</lparam></gate>
<gate>
<ID>478</ID>
<type>DE_TO</type>
<position>61.5,-93.5</position>
<input>
<ID>IN_0</ID>393 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A11</lparam></gate>
<gate>
<ID>479</ID>
<type>DE_TO</type>
<position>-18,-0.5</position>
<input>
<ID>IN_0</ID>719 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Ck1</lparam></gate>
<gate>
<ID>480</ID>
<type>BE_NOR4</type>
<position>73.5,-84.5</position>
<input>
<ID>IN_0</ID>393 </input>
<input>
<ID>IN_1</ID>392 </input>
<input>
<ID>IN_2</ID>391 </input>
<input>
<ID>IN_3</ID>390 </input>
<output>
<ID>OUT</ID>422 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>482</ID>
<type>DE_TO</type>
<position>73.5,-73.5</position>
<input>
<ID>IN_0</ID>422 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z11-8</lparam></gate>
<gate>
<ID>485</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>244.5,-44.5</position>
<input>
<ID>ENABLE_0</ID>398 </input>
<input>
<ID>IN_0</ID>462 </input>
<input>
<ID>IN_1</ID>461 </input>
<input>
<ID>IN_2</ID>460 </input>
<input>
<ID>IN_3</ID>459 </input>
<output>
<ID>OUT_0</ID>458 </output>
<output>
<ID>OUT_1</ID>457 </output>
<output>
<ID>OUT_2</ID>456 </output>
<output>
<ID>OUT_3</ID>455 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>486</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>248,-35</position>
<input>
<ID>ENABLE_0</ID>394 </input>
<input>
<ID>IN_0</ID>466 </input>
<input>
<ID>IN_1</ID>465 </input>
<input>
<ID>IN_2</ID>464 </input>
<input>
<ID>IN_3</ID>463 </input>
<output>
<ID>OUT_0</ID>455 </output>
<output>
<ID>OUT_1</ID>456 </output>
<output>
<ID>OUT_2</ID>457 </output>
<output>
<ID>OUT_3</ID>458 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>487</ID>
<type>DA_FROM</type>
<position>233,-39.5</position>
<input>
<ID>IN_0</ID>459 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A7</lparam></gate>
<gate>
<ID>488</ID>
<type>DA_FROM</type>
<position>232,-43</position>
<input>
<ID>IN_0</ID>460 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A6</lparam></gate>
<gate>
<ID>489</ID>
<type>DA_FROM</type>
<position>231.5,-46.5</position>
<input>
<ID>IN_0</ID>461 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A5</lparam></gate>
<gate>
<ID>490</ID>
<type>DA_FROM</type>
<position>231.5,-50</position>
<input>
<ID>IN_0</ID>462 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A4</lparam></gate>
<gate>
<ID>491</ID>
<type>DA_FROM</type>
<position>297,-27</position>
<input>
<ID>IN_0</ID>463 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>492</ID>
<type>DA_FROM</type>
<position>293,-26.5</position>
<input>
<ID>IN_0</ID>464 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>493</ID>
<type>DA_FROM</type>
<position>289,-26</position>
<input>
<ID>IN_0</ID>465 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>494</ID>
<type>DA_FROM</type>
<position>286,-26</position>
<input>
<ID>IN_0</ID>466 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>495</ID>
<type>DA_FROM</type>
<position>249,-50.5</position>
<input>
<ID>IN_0</ID>467 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>496</ID>
<type>FF_GND</type>
<position>256.5,-50</position>
<output>
<ID>OUT_0</ID>468 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>497</ID>
<type>FF_GND</type>
<position>255.5,-38.5</position>
<output>
<ID>OUT_0</ID>469 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>498</ID>
<type>AE_FULLADDER_4BIT</type>
<position>261,-89.5</position>
<input>
<ID>IN_0</ID>436 </input>
<input>
<ID>IN_1</ID>438 </input>
<input>
<ID>IN_2</ID>439 </input>
<input>
<ID>IN_3</ID>440 </input>
<input>
<ID>IN_B_0</ID>423 </input>
<input>
<ID>IN_B_1</ID>424 </input>
<input>
<ID>IN_B_2</ID>425 </input>
<input>
<ID>IN_B_3</ID>426 </input>
<output>
<ID>OUT_0</ID>446 </output>
<output>
<ID>OUT_1</ID>447 </output>
<output>
<ID>OUT_2</ID>448 </output>
<output>
<ID>OUT_3</ID>449 </output>
<input>
<ID>carry_in</ID>524 </input>
<output>
<ID>carry_out</ID>523 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>499</ID>
<type>AI_XOR2</type>
<position>282,-68</position>
<input>
<ID>IN_0</ID>445 </input>
<input>
<ID>IN_1</ID>431 </input>
<output>
<ID>OUT</ID>423 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>500</ID>
<type>AI_XOR2</type>
<position>275.5,-68</position>
<input>
<ID>IN_0</ID>445 </input>
<input>
<ID>IN_1</ID>432 </input>
<output>
<ID>OUT</ID>424 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>501</ID>
<type>AI_XOR2</type>
<position>270,-68</position>
<input>
<ID>IN_0</ID>445 </input>
<input>
<ID>IN_1</ID>433 </input>
<output>
<ID>OUT</ID>425 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>502</ID>
<type>AI_XOR2</type>
<position>263,-68</position>
<input>
<ID>IN_0</ID>445 </input>
<input>
<ID>IN_1</ID>434 </input>
<output>
<ID>OUT</ID>426 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>503</ID>
<type>DA_FROM</type>
<position>257,-63</position>
<input>
<ID>IN_0</ID>430 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>504</ID>
<type>DA_FROM</type>
<position>250.5,-62.5</position>
<input>
<ID>IN_0</ID>429 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>505</ID>
<type>DA_FROM</type>
<position>245.5,-62.5</position>
<input>
<ID>IN_0</ID>428 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>506</ID>
<type>DA_FROM</type>
<position>239,-62</position>
<input>
<ID>IN_0</ID>427 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>507</ID>
<type>AI_XOR2</type>
<position>258,-69</position>
<input>
<ID>IN_0</ID>444 </input>
<input>
<ID>IN_1</ID>430 </input>
<output>
<ID>OUT</ID>435 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>508</ID>
<type>AI_XOR2</type>
<position>251.5,-69</position>
<input>
<ID>IN_0</ID>444 </input>
<input>
<ID>IN_1</ID>429 </input>
<output>
<ID>OUT</ID>437 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>509</ID>
<type>AI_XOR2</type>
<position>246.5,-69</position>
<input>
<ID>IN_0</ID>444 </input>
<input>
<ID>IN_1</ID>428 </input>
<output>
<ID>OUT</ID>441 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>510</ID>
<type>AI_XOR2</type>
<position>240,-69</position>
<input>
<ID>IN_0</ID>444 </input>
<input>
<ID>IN_1</ID>427 </input>
<output>
<ID>OUT</ID>442 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>511</ID>
<type>AA_REGISTER4</type>
<position>255.5,-45</position>
<input>
<ID>IN_0</ID>458 </input>
<input>
<ID>IN_1</ID>457 </input>
<input>
<ID>IN_2</ID>456 </input>
<input>
<ID>IN_3</ID>455 </input>
<output>
<ID>OUT_0</ID>431 </output>
<output>
<ID>OUT_1</ID>432 </output>
<output>
<ID>OUT_2</ID>433 </output>
<output>
<ID>OUT_3</ID>434 </output>
<input>
<ID>clear</ID>468 </input>
<input>
<ID>clock</ID>467 </input>
<input>
<ID>count_enable</ID>469 </input>
<input>
<ID>count_up</ID>469 </input>
<input>
<ID>load</ID>470 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>512</ID>
<type>AA_AND2</type>
<position>259,-77.5</position>
<input>
<ID>IN_0</ID>443 </input>
<input>
<ID>IN_1</ID>435 </input>
<output>
<ID>OUT</ID>436 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>513</ID>
<type>AA_AND2</type>
<position>252.5,-78</position>
<input>
<ID>IN_0</ID>443 </input>
<input>
<ID>IN_1</ID>437 </input>
<output>
<ID>OUT</ID>438 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>514</ID>
<type>AA_AND2</type>
<position>247.5,-78</position>
<input>
<ID>IN_0</ID>443 </input>
<input>
<ID>IN_1</ID>441 </input>
<output>
<ID>OUT</ID>439 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>515</ID>
<type>AA_AND2</type>
<position>241,-78</position>
<input>
<ID>IN_0</ID>443 </input>
<input>
<ID>IN_1</ID>442 </input>
<output>
<ID>OUT</ID>440 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>516</ID>
<type>AE_SMALL_INVERTER</type>
<position>236.5,-73.5</position>
<input>
<ID>IN_0</ID>471 </input>
<output>
<ID>OUT_0</ID>443 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>519</ID>
<type>AA_AND4</type>
<position>-113.5,-27.5</position>
<input>
<ID>IN_0</ID>624 </input>
<input>
<ID>IN_1</ID>625 </input>
<input>
<ID>IN_2</ID>626 </input>
<input>
<ID>IN_3</ID>627 </input>
<output>
<ID>OUT</ID>630 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>521</ID>
<type>DA_FROM</type>
<position>267.5,-36.5</position>
<input>
<ID>IN_0</ID>470 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LD Acc</lparam></gate>
<gate>
<ID>522</ID>
<type>DA_FROM</type>
<position>227.5,-73.5</position>
<input>
<ID>IN_0</ID>471 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BZero</lparam></gate>
<gate>
<ID>523</ID>
<type>DE_TO</type>
<position>209.5,-98</position>
<input>
<ID>IN_0</ID>446 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A4</lparam></gate>
<gate>
<ID>524</ID>
<type>DE_TO</type>
<position>204,-96.5</position>
<input>
<ID>IN_0</ID>447 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A5</lparam></gate>
<gate>
<ID>525</ID>
<type>DE_TO</type>
<position>210.5,-95</position>
<input>
<ID>IN_0</ID>448 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A6</lparam></gate>
<gate>
<ID>526</ID>
<type>DE_TO</type>
<position>204.5,-93.5</position>
<input>
<ID>IN_0</ID>449 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A7</lparam></gate>
<gate>
<ID>527</ID>
<type>BE_NOR4</type>
<position>216.5,-84.5</position>
<input>
<ID>IN_0</ID>449 </input>
<input>
<ID>IN_1</ID>448 </input>
<input>
<ID>IN_2</ID>447 </input>
<input>
<ID>IN_3</ID>446 </input>
<output>
<ID>OUT</ID>472 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>528</ID>
<type>DE_TO</type>
<position>216.5,-73.5</position>
<input>
<ID>IN_0</ID>472 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z7-4</lparam></gate>
<gate>
<ID>529</ID>
<type>AA_MUX_2x1</type>
<position>-113.5,-20.5</position>
<input>
<ID>IN_0</ID>315 </input>
<input>
<ID>IN_1</ID>630 </input>
<output>
<ID>OUT</ID>629 </output>
<input>
<ID>SEL_0</ID>631 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>531</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>387,-43.5</position>
<input>
<ID>ENABLE_0</ID>450 </input>
<input>
<ID>IN_0</ID>512 </input>
<input>
<ID>IN_1</ID>511 </input>
<input>
<ID>IN_2</ID>510 </input>
<input>
<ID>IN_3</ID>509 </input>
<output>
<ID>OUT_0</ID>508 </output>
<output>
<ID>OUT_1</ID>507 </output>
<output>
<ID>OUT_2</ID>506 </output>
<output>
<ID>OUT_3</ID>505 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>532</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>390.5,-34</position>
<input>
<ID>ENABLE_0</ID>395 </input>
<input>
<ID>IN_0</ID>516 </input>
<input>
<ID>IN_1</ID>515 </input>
<input>
<ID>IN_2</ID>514 </input>
<input>
<ID>IN_3</ID>513 </input>
<output>
<ID>OUT_0</ID>505 </output>
<output>
<ID>OUT_1</ID>506 </output>
<output>
<ID>OUT_2</ID>507 </output>
<output>
<ID>OUT_3</ID>508 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>533</ID>
<type>DA_FROM</type>
<position>380,-42</position>
<input>
<ID>IN_0</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>534</ID>
<type>DA_FROM</type>
<position>375.5,-43</position>
<input>
<ID>IN_0</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>535</ID>
<type>DA_FROM</type>
<position>370,-44</position>
<input>
<ID>IN_0</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>536</ID>
<type>DA_FROM</type>
<position>364,-45</position>
<input>
<ID>IN_0</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>537</ID>
<type>DA_FROM</type>
<position>441.5,-24.5</position>
<input>
<ID>IN_0</ID>513 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>538</ID>
<type>DA_FROM</type>
<position>437,-22</position>
<input>
<ID>IN_0</ID>514 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>539</ID>
<type>DA_FROM</type>
<position>432.5,-22</position>
<input>
<ID>IN_0</ID>515 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>540</ID>
<type>DA_FROM</type>
<position>428.5,-21</position>
<input>
<ID>IN_0</ID>516 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>541</ID>
<type>DA_FROM</type>
<position>391.5,-49.5</position>
<input>
<ID>IN_0</ID>517 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>542</ID>
<type>FF_GND</type>
<position>399,-49</position>
<output>
<ID>OUT_0</ID>518 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>543</ID>
<type>FF_GND</type>
<position>398,-36.5</position>
<output>
<ID>OUT_0</ID>519 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>544</ID>
<type>AE_FULLADDER_4BIT</type>
<position>403.5,-88.5</position>
<input>
<ID>IN_0</ID>486 </input>
<input>
<ID>IN_1</ID>488 </input>
<input>
<ID>IN_2</ID>489 </input>
<input>
<ID>IN_3</ID>490 </input>
<input>
<ID>IN_B_0</ID>473 </input>
<input>
<ID>IN_B_1</ID>474 </input>
<input>
<ID>IN_B_2</ID>475 </input>
<input>
<ID>IN_B_3</ID>476 </input>
<output>
<ID>OUT_0</ID>496 </output>
<output>
<ID>OUT_1</ID>497 </output>
<output>
<ID>OUT_2</ID>498 </output>
<output>
<ID>OUT_3</ID>499 </output>
<input>
<ID>carry_in</ID>500 </input>
<output>
<ID>carry_out</ID>524 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>545</ID>
<type>AI_XOR2</type>
<position>424.5,-67</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>481 </input>
<output>
<ID>OUT</ID>473 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>546</ID>
<type>AI_XOR2</type>
<position>418,-67</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>482 </input>
<output>
<ID>OUT</ID>474 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>547</ID>
<type>AI_XOR2</type>
<position>412.5,-67</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>483 </input>
<output>
<ID>OUT</ID>475 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>548</ID>
<type>AI_XOR2</type>
<position>405.5,-67</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>484 </input>
<output>
<ID>OUT</ID>476 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>549</ID>
<type>DA_FROM</type>
<position>399.5,-60</position>
<input>
<ID>IN_0</ID>480 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>550</ID>
<type>DA_FROM</type>
<position>393,-59.5</position>
<input>
<ID>IN_0</ID>479 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>551</ID>
<type>DA_FROM</type>
<position>388,-59</position>
<input>
<ID>IN_0</ID>478 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>552</ID>
<type>DA_FROM</type>
<position>381.5,-59</position>
<input>
<ID>IN_0</ID>477 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>553</ID>
<type>AI_XOR2</type>
<position>400.5,-68</position>
<input>
<ID>IN_0</ID>494 </input>
<input>
<ID>IN_1</ID>480 </input>
<output>
<ID>OUT</ID>485 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>554</ID>
<type>AI_XOR2</type>
<position>394,-68</position>
<input>
<ID>IN_0</ID>494 </input>
<input>
<ID>IN_1</ID>479 </input>
<output>
<ID>OUT</ID>487 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>555</ID>
<type>AI_XOR2</type>
<position>389,-68</position>
<input>
<ID>IN_0</ID>494 </input>
<input>
<ID>IN_1</ID>478 </input>
<output>
<ID>OUT</ID>491 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>556</ID>
<type>AI_XOR2</type>
<position>382.5,-68</position>
<input>
<ID>IN_0</ID>494 </input>
<input>
<ID>IN_1</ID>477 </input>
<output>
<ID>OUT</ID>492 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>557</ID>
<type>AA_REGISTER4</type>
<position>398,-44</position>
<input>
<ID>IN_0</ID>508 </input>
<input>
<ID>IN_1</ID>507 </input>
<input>
<ID>IN_2</ID>506 </input>
<input>
<ID>IN_3</ID>505 </input>
<output>
<ID>OUT_0</ID>481 </output>
<output>
<ID>OUT_1</ID>482 </output>
<output>
<ID>OUT_2</ID>483 </output>
<output>
<ID>OUT_3</ID>484 </output>
<input>
<ID>clear</ID>518 </input>
<input>
<ID>clock</ID>517 </input>
<input>
<ID>count_enable</ID>519 </input>
<input>
<ID>count_up</ID>519 </input>
<input>
<ID>load</ID>520 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>558</ID>
<type>AA_AND2</type>
<position>401.5,-76.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>485 </input>
<output>
<ID>OUT</ID>486 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>559</ID>
<type>AA_AND2</type>
<position>395,-77</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>487 </input>
<output>
<ID>OUT</ID>488 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>560</ID>
<type>AA_AND2</type>
<position>390,-77</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>491 </input>
<output>
<ID>OUT</ID>489 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>561</ID>
<type>AA_AND2</type>
<position>383.5,-77</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>490 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>562</ID>
<type>AE_SMALL_INVERTER</type>
<position>379,-72.5</position>
<input>
<ID>IN_0</ID>521 </input>
<output>
<ID>OUT_0</ID>493 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>563</ID>
<type>DA_FROM</type>
<position>-122,-20.5</position>
<input>
<ID>IN_0</ID>631 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID StatEn</lparam></gate>
<gate>
<ID>564</ID>
<type>AE_OR2</type>
<position>433.5,-66.5</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>494 </input>
<output>
<ID>OUT</ID>500 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>565</ID>
<type>AA_MUX_2x1</type>
<position>-115.5,-69.5</position>
<input>
<ID>IN_0</ID>303 </input>
<input>
<ID>IN_1</ID>336 </input>
<output>
<ID>OUT</ID>662 </output>
<input>
<ID>SEL_0</ID>632 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>566</ID>
<type>DA_FROM</type>
<position>-124,-69.5</position>
<input>
<ID>IN_0</ID>632 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID StatEn</lparam></gate>
<gate>
<ID>567</ID>
<type>DA_FROM</type>
<position>408,-34.5</position>
<input>
<ID>IN_0</ID>520 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LD Acc</lparam></gate>
<gate>
<ID>568</ID>
<type>DA_FROM</type>
<position>370,-72.5</position>
<input>
<ID>IN_0</ID>521 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BZero</lparam></gate>
<gate>
<ID>569</ID>
<type>DE_TO</type>
<position>352,-97</position>
<input>
<ID>IN_0</ID>496 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>570</ID>
<type>DE_TO</type>
<position>346.5,-95.5</position>
<input>
<ID>IN_0</ID>497 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>571</ID>
<type>DE_TO</type>
<position>353,-94</position>
<input>
<ID>IN_0</ID>498 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>572</ID>
<type>DE_TO</type>
<position>347,-92.5</position>
<input>
<ID>IN_0</ID>499 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>573</ID>
<type>BE_NOR4</type>
<position>359,-83.5</position>
<input>
<ID>IN_0</ID>499 </input>
<input>
<ID>IN_1</ID>498 </input>
<input>
<ID>IN_2</ID>497 </input>
<input>
<ID>IN_3</ID>496 </input>
<output>
<ID>OUT</ID>522 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>574</ID>
<type>DE_TO</type>
<position>359,-72.5</position>
<input>
<ID>IN_0</ID>522 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z3-0</lparam></gate>
<gate>
<ID>575</ID>
<type>AA_MUX_2x1</type>
<position>-101,-84.5</position>
<input>
<ID>IN_0</ID>294 </input>
<input>
<ID>IN_1</ID>692 </input>
<output>
<ID>OUT</ID>669 </output>
<input>
<ID>SEL_0</ID>668 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>576</ID>
<type>DA_FROM</type>
<position>-113,-84.5</position>
<input>
<ID>IN_0</ID>668 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID StatEn</lparam></gate>
<gate>
<ID>577</ID>
<type>AA_MUX_2x1</type>
<position>-79.5,-83.5</position>
<input>
<ID>IN_0</ID>298 </input>
<input>
<ID>IN_1</ID>704 </input>
<output>
<ID>OUT</ID>703 </output>
<input>
<ID>SEL_0</ID>702 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>578</ID>
<type>DA_FROM</type>
<position>-89.5,-69.5</position>
<input>
<ID>IN_0</ID>702 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID StatEn</lparam></gate>
<gate>
<ID>586</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>427,-43.5</position>
<input>
<ID>ENABLE_0</ID>531 </input>
<input>
<ID>IN_0</ID>481 </input>
<input>
<ID>IN_1</ID>482 </input>
<input>
<ID>IN_2</ID>483 </input>
<input>
<ID>IN_3</ID>484 </input>
<output>
<ID>OUT_0</ID>513 </output>
<output>
<ID>OUT_1</ID>514 </output>
<output>
<ID>OUT_2</ID>515 </output>
<output>
<ID>OUT_3</ID>516 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>588</ID>
<type>DA_FROM</type>
<position>423,-39.5</position>
<input>
<ID>IN_0</ID>531 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Acc-Bus</lparam></gate>
<gate>
<ID>589</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>284,-44.5</position>
<input>
<ID>ENABLE_0</ID>532 </input>
<input>
<ID>IN_0</ID>431 </input>
<input>
<ID>IN_1</ID>432 </input>
<input>
<ID>IN_2</ID>433 </input>
<input>
<ID>IN_3</ID>434 </input>
<output>
<ID>OUT_0</ID>463 </output>
<output>
<ID>OUT_1</ID>464 </output>
<output>
<ID>OUT_2</ID>465 </output>
<output>
<ID>OUT_3</ID>466 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>590</ID>
<type>DA_FROM</type>
<position>274,-40</position>
<input>
<ID>IN_0</ID>532 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Acc-Bus</lparam></gate>
<gate>
<ID>591</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>141.5,-44.5</position>
<input>
<ID>ENABLE_0</ID>533 </input>
<input>
<ID>IN_0</ID>375 </input>
<input>
<ID>IN_1</ID>376 </input>
<input>
<ID>IN_2</ID>377 </input>
<input>
<ID>IN_3</ID>378 </input>
<output>
<ID>OUT_0</ID>407 </output>
<output>
<ID>OUT_1</ID>408 </output>
<output>
<ID>OUT_2</ID>409 </output>
<output>
<ID>OUT_3</ID>410 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>592</ID>
<type>DA_FROM</type>
<position>139,-40</position>
<input>
<ID>IN_0</ID>533 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Acc-Bus</lparam></gate>
<gate>
<ID>593</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>-15,-44</position>
<input>
<ID>ENABLE_0</ID>534 </input>
<input>
<ID>IN_0</ID>317 </input>
<input>
<ID>IN_1</ID>318 </input>
<input>
<ID>IN_2</ID>319 </input>
<input>
<ID>IN_3</ID>320 </input>
<output>
<ID>OUT_0</ID>351 </output>
<output>
<ID>OUT_1</ID>352 </output>
<output>
<ID>OUT_2</ID>353 </output>
<output>
<ID>OUT_3</ID>354 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>594</ID>
<type>DA_FROM</type>
<position>-17.5,-39.5</position>
<input>
<ID>IN_0</ID>534 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Acc-Bus</lparam></gate>
<gate>
<ID>596</ID>
<type>DA_FROM</type>
<position>442,-60.5</position>
<input>
<ID>IN_0</ID>495 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBA</lparam></gate>
<gate>
<ID>597</ID>
<type>DA_FROM</type>
<position>440.5,-56</position>
<input>
<ID>IN_0</ID>494 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBB</lparam></gate>
<gate>
<ID>599</ID>
<type>DA_FROM</type>
<position>298,-60.5</position>
<input>
<ID>IN_0</ID>445 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBA</lparam></gate>
<gate>
<ID>600</ID>
<type>DA_FROM</type>
<position>296.5,-56</position>
<input>
<ID>IN_0</ID>444 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBB</lparam></gate>
<gate>
<ID>601</ID>
<type>DA_FROM</type>
<position>147.5,-60.5</position>
<input>
<ID>IN_0</ID>389 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBA</lparam></gate>
<gate>
<ID>602</ID>
<type>DA_FROM</type>
<position>146,-56</position>
<input>
<ID>IN_0</ID>388 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBB</lparam></gate>
<gate>
<ID>603</ID>
<type>DA_FROM</type>
<position>-109,-37.5</position>
<input>
<ID>IN_0</ID>626 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z7-4</lparam></gate>
<gate>
<ID>604</ID>
<type>DA_FROM</type>
<position>-106,-37.5</position>
<input>
<ID>IN_0</ID>627 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Z3-0</lparam></gate>
<gate>
<ID>605</ID>
<type>DA_FROM</type>
<position>-6,-56.5</position>
<input>
<ID>IN_0</ID>332 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBA</lparam></gate>
<gate>
<ID>606</ID>
<type>DA_FROM</type>
<position>-8,-52.5</position>
<input>
<ID>IN_0</ID>331 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SUBB</lparam></gate>
<gate>
<ID>608</ID>
<type>DA_FROM</type>
<position>-57,-38</position>
<input>
<ID>IN_0</ID>537 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD Acc</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_LABEL</type>
<position>4,-10</position>
<gparam>LABEL_TEXT Accumulator</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>660</ID>
<type>AA_TOGGLE</type>
<position>-18,-6.5</position>
<output>
<ID>OUT_0</ID>719 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>335</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-37.5,-89</position>
<input>
<ID>IN_0</ID>322 </input>
<input>
<ID>IN_1</ID>324 </input>
<input>
<ID>IN_2</ID>325 </input>
<input>
<ID>IN_3</ID>326 </input>
<input>
<ID>IN_B_0</ID>287 </input>
<input>
<ID>IN_B_1</ID>288 </input>
<input>
<ID>IN_B_2</ID>289 </input>
<input>
<ID>IN_B_3</ID>290 </input>
<output>
<ID>OUT_0</ID>661 </output>
<output>
<ID>OUT_1</ID>334 </output>
<output>
<ID>OUT_2</ID>335 </output>
<output>
<ID>OUT_3</ID>336 </output>
<input>
<ID>carry_in</ID>414 </input>
<output>
<ID>carry_out</ID>692 </output>
<output>
<ID>overflow</ID>704 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>336</ID>
<type>AE_DFF_LOW</type>
<position>-98,-79</position>
<input>
<ID>IN_0</ID>669 </input>
<output>
<ID>OUT_0</ID>294 </output>
<input>
<ID>clear</ID>292 </input>
<input>
<ID>clock</ID>293 </input>
<input>
<ID>set</ID>291 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>337</ID>
<type>EE_VDD</type>
<position>-104,-79</position>
<output>
<ID>OUT_0</ID>291 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>338</ID>
<type>AI_XOR2</type>
<position>-16.5,-67.5</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>317 </input>
<output>
<ID>OUT</ID>287 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>339</ID>
<type>AI_XOR2</type>
<position>-23,-67.5</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>318 </input>
<output>
<ID>OUT</ID>288 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>340</ID>
<type>AI_XOR2</type>
<position>-28.5,-67.5</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>319 </input>
<output>
<ID>OUT</ID>289 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>341</ID>
<type>AI_XOR2</type>
<position>-35.5,-67.5</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>320 </input>
<output>
<ID>OUT</ID>290 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>342</ID>
<type>EE_VDD</type>
<position>-88,-79</position>
<output>
<ID>OUT_0</ID>292 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>343</ID>
<type>DA_FROM</type>
<position>-41.5,-62</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>344</ID>
<type>DA_FROM</type>
<position>-48,-61</position>
<input>
<ID>IN_0</ID>309 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>345</ID>
<type>DA_FROM</type>
<position>-53,-61.5</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>346</ID>
<type>DA_FROM</type>
<position>-59.5,-59.5</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>347</ID>
<type>GA_LED</type>
<position>-103.5,-90</position>
<input>
<ID>N_in1</ID>704 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>348</ID>
<type>DA_FROM</type>
<position>-97,-84.5</position>
<input>
<ID>IN_0</ID>293 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>349</ID>
<type>GA_LED</type>
<position>-100,-71.5</position>
<input>
<ID>N_in2</ID>294 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>350</ID>
<type>GA_LED</type>
<position>-107,-88</position>
<input>
<ID>N_in1</ID>692 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>351</ID>
<type>AI_XOR2</type>
<position>-40.5,-68.5</position>
<input>
<ID>IN_0</ID>331 </input>
<input>
<ID>IN_1</ID>310 </input>
<output>
<ID>OUT</ID>321 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>352</ID>
<type>AI_XOR2</type>
<position>-47,-68.5</position>
<input>
<ID>IN_0</ID>331 </input>
<input>
<ID>IN_1</ID>309 </input>
<output>
<ID>OUT</ID>323 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>353</ID>
<type>AI_XOR2</type>
<position>-52,-68.5</position>
<input>
<ID>IN_0</ID>331 </input>
<input>
<ID>IN_1</ID>308 </input>
<output>
<ID>OUT</ID>327 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>354</ID>
<type>AI_XOR2</type>
<position>-58.5,-68.5</position>
<input>
<ID>IN_0</ID>331 </input>
<input>
<ID>IN_1</ID>307 </input>
<output>
<ID>OUT</ID>328 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>355</ID>
<type>DE_TO</type>
<position>-103,-74.5</position>
<input>
<ID>IN_0</ID>294 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Carry</lparam></gate>
<gate>
<ID>356</ID>
<type>AE_DFF_LOW</type>
<position>-77.5,-78.5</position>
<input>
<ID>IN_0</ID>703 </input>
<output>
<ID>OUT_0</ID>298 </output>
<input>
<ID>clear</ID>296 </input>
<input>
<ID>clock</ID>297 </input>
<input>
<ID>set</ID>295 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>357</ID>
<type>EE_VDD</type>
<position>-83.5,-78.5</position>
<output>
<ID>OUT_0</ID>295 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>358</ID>
<type>EE_VDD</type>
<position>-70,-78.5</position>
<output>
<ID>OUT_0</ID>296 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>359</ID>
<type>DA_FROM</type>
<position>-76.5,-84</position>
<input>
<ID>IN_0</ID>297 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>360</ID>
<type>GA_LED</type>
<position>-79.5,-71</position>
<input>
<ID>N_in2</ID>298 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>362</ID>
<type>DE_TO</type>
<position>-81.5,-73.5</position>
<input>
<ID>IN_0</ID>298 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID oVerflow</lparam></gate>
<gate>
<ID>364</ID>
<type>AE_DFF_LOW</type>
<position>-109,-60</position>
<input>
<ID>IN_0</ID>662 </input>
<output>
<ID>OUT_0</ID>303 </output>
<input>
<ID>clear</ID>301 </input>
<input>
<ID>clock</ID>302 </input>
<input>
<ID>set</ID>299 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>366</ID>
<type>EE_VDD</type>
<position>-115,-60</position>
<output>
<ID>OUT_0</ID>299 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>368</ID>
<type>EE_VDD</type>
<position>-103,-60</position>
<output>
<ID>OUT_0</ID>301 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>369</ID>
<type>AA_REGISTER4</type>
<position>-43,-44.5</position>
<input>
<ID>IN_0</ID>346 </input>
<input>
<ID>IN_1</ID>345 </input>
<input>
<ID>IN_2</ID>344 </input>
<input>
<ID>IN_3</ID>343 </input>
<output>
<ID>OUT_0</ID>317 </output>
<output>
<ID>OUT_1</ID>318 </output>
<output>
<ID>OUT_2</ID>319 </output>
<output>
<ID>OUT_3</ID>320 </output>
<input>
<ID>clear</ID>356 </input>
<input>
<ID>clock</ID>355 </input>
<input>
<ID>count_enable</ID>357 </input>
<input>
<ID>count_up</ID>357 </input>
<input>
<ID>load</ID>537 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>370</ID>
<type>DA_FROM</type>
<position>-108,-65.5</position>
<input>
<ID>IN_0</ID>302 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>371</ID>
<type>AA_AND2</type>
<position>-39.5,-77</position>
<input>
<ID>IN_0</ID>329 </input>
<input>
<ID>IN_1</ID>321 </input>
<output>
<ID>OUT</ID>322 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>372</ID>
<type>AA_AND2</type>
<position>-46,-77.5</position>
<input>
<ID>IN_0</ID>329 </input>
<input>
<ID>IN_1</ID>323 </input>
<output>
<ID>OUT</ID>324 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>373</ID>
<type>AA_AND2</type>
<position>-51,-77.5</position>
<input>
<ID>IN_0</ID>329 </input>
<input>
<ID>IN_1</ID>327 </input>
<output>
<ID>OUT</ID>325 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>374</ID>
<type>AA_AND2</type>
<position>-57.5,-77.5</position>
<input>
<ID>IN_0</ID>329 </input>
<input>
<ID>IN_1</ID>328 </input>
<output>
<ID>OUT</ID>326 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>375</ID>
<type>GA_LED</type>
<position>-111,-52.5</position>
<input>
<ID>N_in2</ID>303 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>376</ID>
<type>AE_SMALL_INVERTER</type>
<position>-62,-73</position>
<input>
<ID>IN_0</ID>417 </input>
<output>
<ID>OUT_0</ID>329 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>377</ID>
<type>DE_TO</type>
<position>-114,-55.5</position>
<input>
<ID>IN_0</ID>303 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID sigN</lparam></gate>
<gate>
<ID>379</ID>
<type>AE_DFF_LOW</type>
<position>-111.5,-14</position>
<input>
<ID>IN_0</ID>629 </input>
<output>
<ID>OUT_0</ID>315 </output>
<input>
<ID>clear</ID>306 </input>
<input>
<ID>clock</ID>311 </input>
<input>
<ID>set</ID>304 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>381</ID>
<type>EE_VDD</type>
<position>-115.5,-13</position>
<output>
<ID>OUT_0</ID>304 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>382</ID>
<type>DA_FROM</type>
<position>-39,-34.5</position>
<input>
<ID>IN_0</ID>369 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus-Acc</lparam></gate>
<gate>
<ID>383</ID>
<type>EE_VDD</type>
<position>-103.5,-13</position>
<output>
<ID>OUT_0</ID>306 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>384</ID>
<type>DA_FROM</type>
<position>110,-35</position>
<input>
<ID>IN_0</ID>370 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus-Acc</lparam></gate>
<gate>
<ID>385</ID>
<type>DA_FROM</type>
<position>253,-35</position>
<input>
<ID>IN_0</ID>394 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus-Acc</lparam></gate>
<gate>
<ID>386</ID>
<type>DA_FROM</type>
<position>397,-33</position>
<input>
<ID>IN_0</ID>395 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Bus-Acc</lparam></gate>
<gate>
<ID>387</ID>
<type>DA_FROM</type>
<position>-54,-30.5</position>
<input>
<ID>IN_0</ID>396 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Res-Acc</lparam></gate>
<gate>
<ID>388</ID>
<type>DA_FROM</type>
<position>-109,-20.5</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-65,121,-54</points>
<connection>
<GID>435</GID>
<name>IN_0</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-54,140,-54</points>
<intersection>121 0</intersection>
<intersection>128 3</intersection>
<intersection>133.5 7</intersection>
<intersection>140 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128,-65,128,-54</points>
<connection>
<GID>434</GID>
<name>IN_0</name></connection>
<intersection>-54 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>140,-65,140,-54</points>
<connection>
<GID>432</GID>
<name>IN_0</name></connection>
<intersection>-60.5 10</intersection>
<intersection>-54 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>133.5,-65,133.5,-54</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>140,-60.5,145.5,-60.5</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<intersection>140 6</intersection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-98,119.5,-93.5</points>
<connection>
<GID>431</GID>
<name>OUT_0</name></connection>
<intersection>-98 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>68.5,-98,119.5,-98</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>76.5 8</intersection>
<intersection>119.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>76.5,-98,76.5,-87.5</points>
<connection>
<GID>480</GID>
<name>IN_3</name></connection>
<intersection>-98 7</intersection></vsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-96.5,118.5,-93.5</points>
<connection>
<GID>431</GID>
<name>OUT_1</name></connection>
<intersection>-96.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>63,-96.5,118.5,-96.5</points>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<intersection>74.5 8</intersection>
<intersection>118.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>74.5,-96.5,74.5,-87.5</points>
<connection>
<GID>480</GID>
<name>IN_2</name></connection>
<intersection>-96.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-95,117.5,-93.5</points>
<connection>
<GID>431</GID>
<name>OUT_2</name></connection>
<intersection>-95 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>69.5,-95,117.5,-95</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<intersection>72.5 8</intersection>
<intersection>117.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>72.5,-95,72.5,-87.5</points>
<connection>
<GID>480</GID>
<name>IN_1</name></connection>
<intersection>-95 7</intersection></vsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>63.5,-93.5,116.5,-93.5</points>
<connection>
<GID>431</GID>
<name>OUT_3</name></connection>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>70.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>70.5,-93.5,70.5,-87.5</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>-93.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-35,251,-35</points>
<connection>
<GID>486</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>385</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394,-34,394,-33</points>
<intersection>-34 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>393.5,-34,394,-34</points>
<connection>
<GID>532</GID>
<name>ENABLE_0</name></connection>
<intersection>394 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>394,-33,395,-33</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>394 0</intersection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54,-41,-54,-32.5</points>
<connection>
<GID>395</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>387</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-41.5,101.5,-27</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<connection>
<GID>418</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244.5,-41.5,244.5,-33.5</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<connection>
<GID>485</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,-43,108.5,-43</points>
<connection>
<GID>418</GID>
<name>OUT_3</name></connection>
<connection>
<GID>450</GID>
<name>IN_3</name></connection>
<intersection>103.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>103.5,-43,103.5,-37</points>
<connection>
<GID>419</GID>
<name>OUT_0</name></connection>
<intersection>-43 1</intersection></vsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,-44,108.5,-44</points>
<connection>
<GID>418</GID>
<name>OUT_2</name></connection>
<connection>
<GID>450</GID>
<name>IN_2</name></connection>
<intersection>104.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>104.5,-44,104.5,-37</points>
<connection>
<GID>419</GID>
<name>OUT_1</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,-45,108.5,-45</points>
<connection>
<GID>418</GID>
<name>OUT_1</name></connection>
<connection>
<GID>450</GID>
<name>IN_1</name></connection>
<intersection>105.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>105.5,-45,105.5,-37</points>
<connection>
<GID>419</GID>
<name>OUT_2</name></connection>
<intersection>-45 1</intersection></vsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,-46,108.5,-46</points>
<connection>
<GID>418</GID>
<name>OUT_0</name></connection>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<intersection>106.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>106.5,-46,106.5,-37</points>
<connection>
<GID>419</GID>
<name>OUT_3</name></connection>
<intersection>-46 1</intersection></vsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96.5,-43,99.5,-43</points>
<connection>
<GID>418</GID>
<name>IN_3</name></connection>
<connection>
<GID>420</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>92,-44,99.5,-44</points>
<connection>
<GID>418</GID>
<name>IN_2</name></connection>
<connection>
<GID>421</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-45,99.5,-45</points>
<connection>
<GID>418</GID>
<name>IN_1</name></connection>
<connection>
<GID>422</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80.5,-46,99.5,-46</points>
<connection>
<GID>418</GID>
<name>IN_0</name></connection>
<connection>
<GID>423</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-33,106.5,-32.5</points>
<connection>
<GID>419</GID>
<name>IN_3</name></connection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>106.5,-32.5,156,-32.5</points>
<intersection>106.5 0</intersection>
<intersection>156 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>156,-46,156,-27</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>-46 5</intersection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>143.5,-46,156,-46</points>
<connection>
<GID>591</GID>
<name>OUT_0</name></connection>
<intersection>156 3</intersection></hsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,-45,152,-26.5</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<intersection>-45 10</intersection>
<intersection>-31.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>105.5,-31.5,152,-31.5</points>
<intersection>105.5 8</intersection>
<intersection>152 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>105.5,-33,105.5,-31.5</points>
<connection>
<GID>419</GID>
<name>IN_2</name></connection>
<intersection>-31.5 7</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>143.5,-45,152,-45</points>
<connection>
<GID>591</GID>
<name>OUT_1</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-33,104.5,-30</points>
<connection>
<GID>419</GID>
<name>IN_1</name></connection>
<intersection>-30 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-30,148,-30</points>
<intersection>104.5 0</intersection>
<intersection>148 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>148,-44,148,-26</points>
<connection>
<GID>426</GID>
<name>IN_0</name></connection>
<intersection>-44 9</intersection>
<intersection>-30 3</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>143.5,-44,148,-44</points>
<connection>
<GID>591</GID>
<name>OUT_2</name></connection>
<intersection>148 7</intersection></hsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-33,103.5,-28.5</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>-28.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>145,-43,145,-26</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<intersection>-43 4</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-28.5,145,-28.5</points>
<intersection>103.5 0</intersection>
<intersection>145 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>143.5,-43,145,-43</points>
<connection>
<GID>591</GID>
<name>OUT_3</name></connection>
<intersection>145 1</intersection></hsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-50.5,111.5,-49</points>
<connection>
<GID>450</GID>
<name>clock</name></connection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-50.5,111.5,-50.5</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-49,113.5,-49</points>
<connection>
<GID>429</GID>
<name>OUT_0</name></connection>
<connection>
<GID>450</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-40,112.5,-38.5</points>
<connection>
<GID>430</GID>
<name>OUT_0</name></connection>
<connection>
<GID>450</GID>
<name>count_enable</name></connection>
<intersection>-39.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>112.5,-39.5,113.5,-39.5</points>
<intersection>112.5 0</intersection>
<intersection>113.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>113.5,-40,113.5,-39.5</points>
<connection>
<GID>450</GID>
<name>count_up</name></connection>
<intersection>-39.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-29.5,-88.5,110,-88.5</points>
<connection>
<GID>431</GID>
<name>carry_out</name></connection>
<intersection>-29.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-29.5,-88.5,-29.5,-88</points>
<connection>
<GID>335</GID>
<name>carry_in</name></connection>
<intersection>-88.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-40,111.5,-36</points>
<connection>
<GID>450</GID>
<name>load</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,-36,120.5,-36</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-73.5,91.5,-73.5</points>
<connection>
<GID>455</GID>
<name>IN_0</name></connection>
<connection>
<GID>464</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-66.5,-69.5,-64,-69.5</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>-64 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-64,-73,-64,-69.5</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>-69.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88.5,-80.5,-88.5,-64</points>
<connection>
<GID>397</GID>
<name>OUT</name></connection>
<connection>
<GID>467</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-80.5,73.5,-75.5</points>
<connection>
<GID>480</GID>
<name>OUT</name></connection>
<connection>
<GID>482</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-85.5,282,-71</points>
<connection>
<GID>499</GID>
<name>OUT</name></connection>
<intersection>-85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,-85.5,282,-85.5</points>
<connection>
<GID>498</GID>
<name>IN_B_0</name></connection>
<intersection>282 0</intersection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275.5,-84.5,275.5,-71</points>
<connection>
<GID>500</GID>
<name>OUT</name></connection>
<intersection>-84.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>265,-84.5,275.5,-84.5</points>
<intersection>265 4</intersection>
<intersection>275.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>265,-85.5,265,-84.5</points>
<connection>
<GID>498</GID>
<name>IN_B_1</name></connection>
<intersection>-84.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264,-85.5,264,-83.5</points>
<connection>
<GID>498</GID>
<name>IN_B_2</name></connection>
<intersection>-83.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>270,-83.5,270,-71</points>
<connection>
<GID>501</GID>
<name>OUT</name></connection>
<intersection>-83.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>264,-83.5,270,-83.5</points>
<intersection>264 0</intersection>
<intersection>270 1</intersection></hsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263,-85.5,263,-71</points>
<connection>
<GID>498</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>502</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>239,-66,239,-64</points>
<connection>
<GID>506</GID>
<name>IN_0</name></connection>
<connection>
<GID>510</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-66,245.5,-64.5</points>
<connection>
<GID>505</GID>
<name>IN_0</name></connection>
<connection>
<GID>509</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-66,250.5,-64.5</points>
<connection>
<GID>504</GID>
<name>IN_0</name></connection>
<connection>
<GID>508</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257,-66,257,-65</points>
<connection>
<GID>503</GID>
<name>IN_0</name></connection>
<connection>
<GID>507</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-65,281,-46</points>
<connection>
<GID>499</GID>
<name>IN_1</name></connection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259.5,-46,282,-46</points>
<connection>
<GID>511</GID>
<name>OUT_0</name></connection>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274.5,-65,274.5,-45</points>
<connection>
<GID>500</GID>
<name>IN_1</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259.5,-45,282,-45</points>
<connection>
<GID>511</GID>
<name>OUT_1</name></connection>
<connection>
<GID>589</GID>
<name>IN_1</name></connection>
<intersection>274.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269,-65,269,-44</points>
<connection>
<GID>501</GID>
<name>IN_1</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259.5,-44,282,-44</points>
<connection>
<GID>511</GID>
<name>OUT_2</name></connection>
<connection>
<GID>589</GID>
<name>IN_2</name></connection>
<intersection>269 0</intersection></hsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262,-65,262,-43</points>
<connection>
<GID>502</GID>
<name>IN_1</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259.5,-43,282,-43</points>
<connection>
<GID>511</GID>
<name>OUT_3</name></connection>
<connection>
<GID>589</GID>
<name>IN_3</name></connection>
<intersection>262 0</intersection></hsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258,-74.5,258,-72</points>
<connection>
<GID>507</GID>
<name>OUT</name></connection>
<connection>
<GID>512</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259,-85.5,259,-80.5</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<connection>
<GID>512</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251.5,-75,251.5,-72</points>
<connection>
<GID>508</GID>
<name>OUT</name></connection>
<connection>
<GID>513</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258,-85.5,258,-82</points>
<connection>
<GID>498</GID>
<name>IN_1</name></connection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>252.5,-82,258,-82</points>
<intersection>252.5 3</intersection>
<intersection>258 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>252.5,-82,252.5,-81</points>
<connection>
<GID>513</GID>
<name>OUT</name></connection>
<intersection>-82 2</intersection></vsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257,-85.5,257,-83</points>
<connection>
<GID>498</GID>
<name>IN_2</name></connection>
<intersection>-83 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>247.5,-83,247.5,-81</points>
<connection>
<GID>514</GID>
<name>OUT</name></connection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>247.5,-83,257,-83</points>
<intersection>247.5 1</intersection>
<intersection>257 0</intersection></hsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>241,-84,256,-84</points>
<intersection>241 5</intersection>
<intersection>256 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>256,-85.5,256,-84</points>
<connection>
<GID>498</GID>
<name>IN_3</name></connection>
<intersection>-84 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>241,-84,241,-81</points>
<connection>
<GID>515</GID>
<name>OUT</name></connection>
<intersection>-84 2</intersection></vsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246.5,-75,246.5,-72</points>
<connection>
<GID>509</GID>
<name>OUT</name></connection>
<connection>
<GID>514</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-75,240,-72</points>
<connection>
<GID>510</GID>
<name>OUT</name></connection>
<connection>
<GID>515</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-75,242,-73.5</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>238.5,-73.5,260,-73.5</points>
<connection>
<GID>516</GID>
<name>OUT_0</name></connection>
<intersection>242 0</intersection>
<intersection>248.5 3</intersection>
<intersection>253.5 5</intersection>
<intersection>260 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>248.5,-75,248.5,-73.5</points>
<connection>
<GID>514</GID>
<name>IN_0</name></connection>
<intersection>-73.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>253.5,-75,253.5,-73.5</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<intersection>-73.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>260,-74.5,260,-73.5</points>
<connection>
<GID>512</GID>
<name>IN_0</name></connection>
<intersection>-73.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241,-66,241,-55</points>
<connection>
<GID>510</GID>
<name>IN_0</name></connection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241,-55,259,-55</points>
<intersection>241 0</intersection>
<intersection>247.5 7</intersection>
<intersection>252.5 6</intersection>
<intersection>259 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>259,-66,259,-55</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<intersection>-56 10</intersection>
<intersection>-55 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>252.5,-66,252.5,-55</points>
<connection>
<GID>508</GID>
<name>IN_0</name></connection>
<intersection>-55 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>247.5,-66,247.5,-55</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>259,-56,294.5,-56</points>
<connection>
<GID>600</GID>
<name>IN_0</name></connection>
<intersection>259 5</intersection></hsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264,-65,264,-54</points>
<connection>
<GID>502</GID>
<name>IN_0</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264,-54,283,-54</points>
<intersection>264 0</intersection>
<intersection>271 3</intersection>
<intersection>276.5 7</intersection>
<intersection>283 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>271,-65,271,-54</points>
<connection>
<GID>501</GID>
<name>IN_0</name></connection>
<intersection>-54 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>283,-65,283,-54</points>
<connection>
<GID>499</GID>
<name>IN_0</name></connection>
<intersection>-60.5 10</intersection>
<intersection>-54 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>276.5,-65,276.5,-54</points>
<connection>
<GID>500</GID>
<name>IN_0</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>283,-60.5,296,-60.5</points>
<connection>
<GID>599</GID>
<name>IN_0</name></connection>
<intersection>283 6</intersection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262.5,-98,262.5,-93.5</points>
<connection>
<GID>498</GID>
<name>OUT_0</name></connection>
<intersection>-98 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>211.5,-98,262.5,-98</points>
<connection>
<GID>523</GID>
<name>IN_0</name></connection>
<intersection>219.5 8</intersection>
<intersection>262.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>219.5,-98,219.5,-87.5</points>
<connection>
<GID>527</GID>
<name>IN_3</name></connection>
<intersection>-98 7</intersection></vsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,-96.5,261.5,-93.5</points>
<connection>
<GID>498</GID>
<name>OUT_1</name></connection>
<intersection>-96.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>206,-96.5,261.5,-96.5</points>
<connection>
<GID>524</GID>
<name>IN_0</name></connection>
<intersection>217.5 8</intersection>
<intersection>261.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>217.5,-96.5,217.5,-87.5</points>
<connection>
<GID>527</GID>
<name>IN_2</name></connection>
<intersection>-96.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260.5,-95,260.5,-93.5</points>
<connection>
<GID>498</GID>
<name>OUT_2</name></connection>
<intersection>-95 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>212.5,-95,260.5,-95</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<intersection>215.5 8</intersection>
<intersection>260.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>215.5,-95,215.5,-87.5</points>
<connection>
<GID>527</GID>
<name>IN_1</name></connection>
<intersection>-95 7</intersection></vsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>206.5,-93.5,259.5,-93.5</points>
<connection>
<GID>498</GID>
<name>OUT_3</name></connection>
<connection>
<GID>526</GID>
<name>IN_0</name></connection>
<intersection>213.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>213.5,-93.5,213.5,-87.5</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<intersection>-93.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>387,-40.5,387,-30.5</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<connection>
<GID>531</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>246.5,-43,251.5,-43</points>
<connection>
<GID>485</GID>
<name>OUT_3</name></connection>
<connection>
<GID>511</GID>
<name>IN_3</name></connection>
<intersection>246.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>246.5,-43,246.5,-37</points>
<connection>
<GID>486</GID>
<name>OUT_0</name></connection>
<intersection>-43 1</intersection></vsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>246.5,-44,251.5,-44</points>
<connection>
<GID>485</GID>
<name>OUT_2</name></connection>
<connection>
<GID>511</GID>
<name>IN_2</name></connection>
<intersection>247.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>247.5,-44,247.5,-37</points>
<connection>
<GID>486</GID>
<name>OUT_1</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>246.5,-45,251.5,-45</points>
<connection>
<GID>485</GID>
<name>OUT_1</name></connection>
<connection>
<GID>511</GID>
<name>IN_1</name></connection>
<intersection>248.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>248.5,-45,248.5,-37</points>
<connection>
<GID>486</GID>
<name>OUT_2</name></connection>
<intersection>-45 1</intersection></vsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>246.5,-46,251.5,-46</points>
<connection>
<GID>485</GID>
<name>OUT_0</name></connection>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<intersection>249.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>249.5,-46,249.5,-37</points>
<connection>
<GID>486</GID>
<name>OUT_3</name></connection>
<intersection>-46 1</intersection></vsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235,-39.5,242.5,-39.5</points>
<connection>
<GID>487</GID>
<name>IN_0</name></connection>
<intersection>242.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>242.5,-43,242.5,-39.5</points>
<connection>
<GID>485</GID>
<name>IN_3</name></connection>
<intersection>-39.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>234,-44,242.5,-44</points>
<connection>
<GID>485</GID>
<name>IN_2</name></connection>
<intersection>234 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>234,-44,234,-43</points>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<intersection>-44 0</intersection></vsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>233.5,-45,242.5,-45</points>
<connection>
<GID>485</GID>
<name>IN_1</name></connection>
<intersection>233.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>233.5,-46.5,233.5,-45</points>
<connection>
<GID>489</GID>
<name>IN_0</name></connection>
<intersection>-45 1</intersection></vsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>233.5,-50,242.5,-50</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<intersection>242.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>242.5,-50,242.5,-46</points>
<connection>
<GID>485</GID>
<name>IN_0</name></connection>
<intersection>-50 1</intersection></vsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,-33,249.5,-32</points>
<connection>
<GID>486</GID>
<name>IN_3</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>249.5,-32,297,-32</points>
<intersection>249.5 0</intersection>
<intersection>297 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>297,-46,297,-29</points>
<connection>
<GID>491</GID>
<name>IN_0</name></connection>
<intersection>-46 5</intersection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>286,-46,297,-46</points>
<connection>
<GID>589</GID>
<name>OUT_0</name></connection>
<intersection>297 3</intersection></hsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-45,293,-28.5</points>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<intersection>-45 10</intersection>
<intersection>-31 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>248.5,-31,293,-31</points>
<intersection>248.5 8</intersection>
<intersection>293 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>248.5,-33,248.5,-31</points>
<connection>
<GID>486</GID>
<name>IN_2</name></connection>
<intersection>-31 7</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>286,-45,293,-45</points>
<connection>
<GID>589</GID>
<name>OUT_1</name></connection>
<intersection>293 0</intersection></hsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247.5,-33,247.5,-30</points>
<connection>
<GID>486</GID>
<name>IN_1</name></connection>
<intersection>-30 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>247.5,-30,289,-30</points>
<intersection>247.5 0</intersection>
<intersection>289 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>289,-44,289,-28</points>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<intersection>-44 9</intersection>
<intersection>-30 3</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>286,-44,289,-44</points>
<connection>
<GID>589</GID>
<name>OUT_2</name></connection>
<intersection>289 7</intersection></hsegment></shape></wire>
<wire>
<ID>466</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246.5,-33,246.5,-29</points>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<intersection>-29 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>286,-43,286,-28</points>
<connection>
<GID>589</GID>
<name>OUT_3</name></connection>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>246.5,-29,286,-29</points>
<intersection>246.5 0</intersection>
<intersection>286 1</intersection></hsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>254.5,-50.5,254.5,-49</points>
<connection>
<GID>511</GID>
<name>clock</name></connection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>251,-50.5,254.5,-50.5</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>254.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256.5,-49,256.5,-49</points>
<connection>
<GID>496</GID>
<name>OUT_0</name></connection>
<connection>
<GID>511</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>469</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>255.5,-40,256.5,-40</points>
<connection>
<GID>511</GID>
<name>count_up</name></connection>
<connection>
<GID>511</GID>
<name>count_enable</name></connection>
<intersection>255.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>255.5,-40,255.5,-39.5</points>
<connection>
<GID>497</GID>
<name>OUT_0</name></connection>
<intersection>-40 3</intersection></vsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>254.5,-40,254.5,-36.5</points>
<connection>
<GID>511</GID>
<name>load</name></connection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>254.5,-36.5,265.5,-36.5</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<intersection>254.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>229.5,-73.5,234.5,-73.5</points>
<connection>
<GID>516</GID>
<name>IN_0</name></connection>
<connection>
<GID>522</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216.5,-80.5,216.5,-75.5</points>
<connection>
<GID>527</GID>
<name>OUT</name></connection>
<connection>
<GID>528</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>424.5,-84.5,424.5,-70</points>
<connection>
<GID>545</GID>
<name>OUT</name></connection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408.5,-84.5,424.5,-84.5</points>
<connection>
<GID>544</GID>
<name>IN_B_0</name></connection>
<intersection>424.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>418,-83.5,418,-70</points>
<connection>
<GID>546</GID>
<name>OUT</name></connection>
<intersection>-83.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>407.5,-83.5,418,-83.5</points>
<intersection>407.5 4</intersection>
<intersection>418 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>407.5,-84.5,407.5,-83.5</points>
<connection>
<GID>544</GID>
<name>IN_B_1</name></connection>
<intersection>-83.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>406.5,-84.5,406.5,-82.5</points>
<connection>
<GID>544</GID>
<name>IN_B_2</name></connection>
<intersection>-82.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>412.5,-82.5,412.5,-70</points>
<connection>
<GID>547</GID>
<name>OUT</name></connection>
<intersection>-82.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>406.5,-82.5,412.5,-82.5</points>
<intersection>406.5 0</intersection>
<intersection>412.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>405.5,-84.5,405.5,-70</points>
<connection>
<GID>544</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>548</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>381.5,-65,381.5,-61</points>
<connection>
<GID>552</GID>
<name>IN_0</name></connection>
<connection>
<GID>556</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>388,-65,388,-61</points>
<connection>
<GID>551</GID>
<name>IN_0</name></connection>
<connection>
<GID>555</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393,-65,393,-61.5</points>
<connection>
<GID>550</GID>
<name>IN_0</name></connection>
<connection>
<GID>554</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>399.5,-65,399.5,-62</points>
<connection>
<GID>549</GID>
<name>IN_0</name></connection>
<connection>
<GID>553</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>423.5,-64,423.5,-45</points>
<connection>
<GID>545</GID>
<name>IN_1</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>402,-45,425,-45</points>
<connection>
<GID>557</GID>
<name>OUT_0</name></connection>
<connection>
<GID>586</GID>
<name>IN_0</name></connection>
<intersection>423.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>417,-64,417,-44</points>
<connection>
<GID>546</GID>
<name>IN_1</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>402,-44,425,-44</points>
<connection>
<GID>557</GID>
<name>OUT_1</name></connection>
<connection>
<GID>586</GID>
<name>IN_1</name></connection>
<intersection>417 0</intersection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>411.5,-64,411.5,-43</points>
<connection>
<GID>547</GID>
<name>IN_1</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>402,-43,425,-43</points>
<connection>
<GID>557</GID>
<name>OUT_2</name></connection>
<connection>
<GID>586</GID>
<name>IN_2</name></connection>
<intersection>411.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>404.5,-64,404.5,-42</points>
<connection>
<GID>548</GID>
<name>IN_1</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>402,-42,425,-42</points>
<connection>
<GID>557</GID>
<name>OUT_3</name></connection>
<connection>
<GID>586</GID>
<name>IN_3</name></connection>
<intersection>404.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400.5,-73.5,400.5,-71</points>
<connection>
<GID>553</GID>
<name>OUT</name></connection>
<connection>
<GID>558</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>401.5,-84.5,401.5,-79.5</points>
<connection>
<GID>544</GID>
<name>IN_0</name></connection>
<connection>
<GID>558</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>394,-74,394,-71</points>
<connection>
<GID>554</GID>
<name>OUT</name></connection>
<connection>
<GID>559</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400.5,-84.5,400.5,-81</points>
<connection>
<GID>544</GID>
<name>IN_1</name></connection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>395,-81,400.5,-81</points>
<intersection>395 3</intersection>
<intersection>400.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>395,-81,395,-80</points>
<connection>
<GID>559</GID>
<name>OUT</name></connection>
<intersection>-81 2</intersection></vsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>399.5,-84.5,399.5,-82</points>
<connection>
<GID>544</GID>
<name>IN_2</name></connection>
<intersection>-82 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>390,-82,390,-80</points>
<connection>
<GID>560</GID>
<name>OUT</name></connection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>390,-82,399.5,-82</points>
<intersection>390 1</intersection>
<intersection>399.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398.5,-84.5,398.5,-83</points>
<connection>
<GID>544</GID>
<name>IN_3</name></connection>
<intersection>-83 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>383.5,-83,383.5,-80</points>
<connection>
<GID>561</GID>
<name>OUT</name></connection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>383.5,-83,398.5,-83</points>
<intersection>383.5 1</intersection>
<intersection>398.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>389,-74,389,-71</points>
<connection>
<GID>555</GID>
<name>OUT</name></connection>
<connection>
<GID>560</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>382.5,-74,382.5,-71</points>
<connection>
<GID>556</GID>
<name>OUT</name></connection>
<connection>
<GID>561</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384.5,-74,384.5,-72.5</points>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381,-72.5,402.5,-72.5</points>
<connection>
<GID>562</GID>
<name>OUT_0</name></connection>
<intersection>384.5 0</intersection>
<intersection>391 3</intersection>
<intersection>396 5</intersection>
<intersection>402.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>391,-74,391,-72.5</points>
<connection>
<GID>560</GID>
<name>IN_0</name></connection>
<intersection>-72.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>396,-74,396,-72.5</points>
<connection>
<GID>559</GID>
<name>IN_0</name></connection>
<intersection>-72.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>402.5,-73.5,402.5,-72.5</points>
<connection>
<GID>558</GID>
<name>IN_0</name></connection>
<intersection>-72.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>383.5,-65,383.5,-54</points>
<connection>
<GID>556</GID>
<name>IN_0</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>383.5,-54,432.5,-54</points>
<intersection>383.5 0</intersection>
<intersection>390 7</intersection>
<intersection>395 6</intersection>
<intersection>401.5 5</intersection>
<intersection>432.5 9</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>401.5,-65,401.5,-54</points>
<connection>
<GID>553</GID>
<name>IN_0</name></connection>
<intersection>-54 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>395,-65,395,-54</points>
<connection>
<GID>554</GID>
<name>IN_0</name></connection>
<intersection>-54 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>390,-65,390,-54</points>
<connection>
<GID>555</GID>
<name>IN_0</name></connection>
<intersection>-54 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>432.5,-63.5,432.5,-54</points>
<connection>
<GID>564</GID>
<name>IN_1</name></connection>
<intersection>-56 10</intersection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>432.5,-56,438.5,-56</points>
<connection>
<GID>597</GID>
<name>IN_0</name></connection>
<intersection>432.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>406.5,-64,406.5,-53</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>406.5,-53,434.5,-53</points>
<intersection>406.5 0</intersection>
<intersection>413.5 3</intersection>
<intersection>419 7</intersection>
<intersection>425.5 6</intersection>
<intersection>434.5 9</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>413.5,-64,413.5,-53</points>
<connection>
<GID>547</GID>
<name>IN_0</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>425.5,-64,425.5,-53</points>
<connection>
<GID>545</GID>
<name>IN_0</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>419,-64,419,-53</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>434.5,-63.5,434.5,-53</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<intersection>-60.5 10</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>434.5,-60.5,440,-60.5</points>
<connection>
<GID>596</GID>
<name>IN_0</name></connection>
<intersection>434.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>405,-97,405,-92.5</points>
<connection>
<GID>544</GID>
<name>OUT_0</name></connection>
<intersection>-97 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>354,-97,405,-97</points>
<connection>
<GID>569</GID>
<name>IN_0</name></connection>
<intersection>362 8</intersection>
<intersection>405 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>362,-97,362,-86.5</points>
<connection>
<GID>573</GID>
<name>IN_3</name></connection>
<intersection>-97 7</intersection></vsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>404,-95.5,404,-92.5</points>
<connection>
<GID>544</GID>
<name>OUT_1</name></connection>
<intersection>-95.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>348.5,-95.5,404,-95.5</points>
<connection>
<GID>570</GID>
<name>IN_0</name></connection>
<intersection>360 8</intersection>
<intersection>404 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>360,-95.5,360,-86.5</points>
<connection>
<GID>573</GID>
<name>IN_2</name></connection>
<intersection>-95.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>403,-94,403,-92.5</points>
<connection>
<GID>544</GID>
<name>OUT_2</name></connection>
<intersection>-94 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>355,-94,403,-94</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>358 8</intersection>
<intersection>403 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>358,-94,358,-86.5</points>
<connection>
<GID>573</GID>
<name>IN_1</name></connection>
<intersection>-94 7</intersection></vsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>349,-92.5,402,-92.5</points>
<connection>
<GID>544</GID>
<name>OUT_3</name></connection>
<connection>
<GID>572</GID>
<name>IN_0</name></connection>
<intersection>356 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>356,-92.5,356,-86.5</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<intersection>-92.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>433.5,-87.5,433.5,-69.5</points>
<connection>
<GID>564</GID>
<name>OUT</name></connection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>411.5,-87.5,433.5,-87.5</points>
<connection>
<GID>544</GID>
<name>carry_in</name></connection>
<intersection>433.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>389,-42,394,-42</points>
<connection>
<GID>531</GID>
<name>OUT_3</name></connection>
<connection>
<GID>557</GID>
<name>IN_3</name></connection>
<intersection>389 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>389,-42,389,-36</points>
<connection>
<GID>532</GID>
<name>OUT_0</name></connection>
<intersection>-42 1</intersection></vsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>389,-43,394,-43</points>
<connection>
<GID>531</GID>
<name>OUT_2</name></connection>
<connection>
<GID>557</GID>
<name>IN_2</name></connection>
<intersection>390 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>390,-43,390,-36</points>
<connection>
<GID>532</GID>
<name>OUT_1</name></connection>
<intersection>-43 1</intersection></vsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>389,-44,394,-44</points>
<connection>
<GID>531</GID>
<name>OUT_1</name></connection>
<connection>
<GID>557</GID>
<name>IN_1</name></connection>
<intersection>391 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>391,-44,391,-36</points>
<connection>
<GID>532</GID>
<name>OUT_2</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>389,-45,394,-45</points>
<connection>
<GID>531</GID>
<name>OUT_0</name></connection>
<connection>
<GID>557</GID>
<name>IN_0</name></connection>
<intersection>392 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>392,-45,392,-36</points>
<connection>
<GID>532</GID>
<name>OUT_3</name></connection>
<intersection>-45 1</intersection></vsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382,-42,385,-42</points>
<connection>
<GID>531</GID>
<name>IN_3</name></connection>
<connection>
<GID>533</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>377.5,-43,385,-43</points>
<connection>
<GID>531</GID>
<name>IN_2</name></connection>
<connection>
<GID>534</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>372,-44,385,-44</points>
<connection>
<GID>531</GID>
<name>IN_1</name></connection>
<connection>
<GID>535</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>366,-45,385,-45</points>
<connection>
<GID>531</GID>
<name>IN_0</name></connection>
<connection>
<GID>536</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>392,-32,392,-31</points>
<connection>
<GID>532</GID>
<name>IN_3</name></connection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>392,-31,441.5,-31</points>
<intersection>392 0</intersection>
<intersection>434.5 4</intersection>
<intersection>441.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>441.5,-31,441.5,-26.5</points>
<connection>
<GID>537</GID>
<name>IN_0</name></connection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>434.5,-45,434.5,-31</points>
<intersection>-45 5</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>429,-45,434.5,-45</points>
<connection>
<GID>586</GID>
<name>OUT_0</name></connection>
<intersection>434.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>437,-30,437,-24</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<intersection>-30 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>391,-30,437,-30</points>
<intersection>391 8</intersection>
<intersection>432 9</intersection>
<intersection>437 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>391,-32,391,-30</points>
<connection>
<GID>532</GID>
<name>IN_2</name></connection>
<intersection>-30 7</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>432,-44,432,-30</points>
<intersection>-44 10</intersection>
<intersection>-30 7</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>429,-44,432,-44</points>
<connection>
<GID>586</GID>
<name>OUT_1</name></connection>
<intersection>432 9</intersection></hsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>390,-32,390,-29</points>
<connection>
<GID>532</GID>
<name>IN_1</name></connection>
<intersection>-29 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>390,-29,432.5,-29</points>
<intersection>390 0</intersection>
<intersection>430.5 8</intersection>
<intersection>432.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>432.5,-29,432.5,-24</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<intersection>-29 3</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>430.5,-43,430.5,-29</points>
<intersection>-43 9</intersection>
<intersection>-29 3</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>429,-43,430.5,-43</points>
<connection>
<GID>586</GID>
<name>OUT_2</name></connection>
<intersection>430.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>389,-32,389,-27.5</points>
<connection>
<GID>532</GID>
<name>IN_0</name></connection>
<intersection>-27.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>428.5,-42,428.5,-23</points>
<connection>
<GID>540</GID>
<name>IN_0</name></connection>
<intersection>-42 3</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>389,-27.5,428.5,-27.5</points>
<intersection>389 0</intersection>
<intersection>428.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>428.5,-42,429,-42</points>
<connection>
<GID>586</GID>
<name>OUT_3</name></connection>
<intersection>428.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397,-49.5,397,-48</points>
<connection>
<GID>557</GID>
<name>clock</name></connection>
<intersection>-49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>393.5,-49.5,397,-49.5</points>
<connection>
<GID>541</GID>
<name>IN_0</name></connection>
<intersection>397 0</intersection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>399,-48,399,-48</points>
<connection>
<GID>542</GID>
<name>OUT_0</name></connection>
<connection>
<GID>557</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398,-39,398,-37.5</points>
<connection>
<GID>543</GID>
<name>OUT_0</name></connection>
<connection>
<GID>557</GID>
<name>count_enable</name></connection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>398,-38.5,399,-38.5</points>
<intersection>398 0</intersection>
<intersection>399 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>399,-39,399,-38.5</points>
<connection>
<GID>557</GID>
<name>count_up</name></connection>
<intersection>-38.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397,-39,397,-34.5</points>
<connection>
<GID>557</GID>
<name>load</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>397,-34.5,406,-34.5</points>
<connection>
<GID>567</GID>
<name>IN_0</name></connection>
<intersection>397 0</intersection></hsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>372,-72.5,377,-72.5</points>
<connection>
<GID>562</GID>
<name>IN_0</name></connection>
<connection>
<GID>568</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>359,-79.5,359,-74.5</points>
<connection>
<GID>573</GID>
<name>OUT</name></connection>
<connection>
<GID>574</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-88.5,253,-88.5</points>
<connection>
<GID>498</GID>
<name>carry_out</name></connection>
<connection>
<GID>431</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>269,-88.5,395.5,-88.5</points>
<connection>
<GID>498</GID>
<name>carry_in</name></connection>
<intersection>395.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>395.5,-88.5,395.5,-87.5</points>
<connection>
<GID>544</GID>
<name>carry_out</name></connection>
<intersection>-88.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427,-40.5,427,-39.5</points>
<connection>
<GID>586</GID>
<name>ENABLE_0</name></connection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425,-39.5,427,-39.5</points>
<connection>
<GID>588</GID>
<name>IN_0</name></connection>
<intersection>427 0</intersection></hsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-41.5,284,-40</points>
<connection>
<GID>589</GID>
<name>ENABLE_0</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-40,284,-40</points>
<connection>
<GID>590</GID>
<name>IN_0</name></connection>
<intersection>284 0</intersection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-41.5,141.5,-40</points>
<connection>
<GID>591</GID>
<name>ENABLE_0</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141,-40,141.5,-40</points>
<connection>
<GID>592</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,-41,-15,-39.5</points>
<connection>
<GID>593</GID>
<name>ENABLE_0</name></connection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15.5,-39.5,-15,-39.5</points>
<connection>
<GID>594</GID>
<name>IN_0</name></connection>
<intersection>-15 0</intersection></hsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-39.5,-44,-38</points>
<connection>
<GID>369</GID>
<name>load</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,-38,-44,-38</points>
<connection>
<GID>608</GID>
<name>IN_0</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-116.5,-35,-116.5,-30.5</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<connection>
<GID>519</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-113.5,-35,-113.5,-33</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<intersection>-33 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-114.5,-33,-114.5,-30.5</points>
<connection>
<GID>519</GID>
<name>IN_1</name></connection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-114.5,-33,-113.5,-33</points>
<intersection>-114.5 1</intersection>
<intersection>-113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-109,-35.5,-109,-33</points>
<connection>
<GID>603</GID>
<name>IN_0</name></connection>
<intersection>-33 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-112.5,-33,-112.5,-30.5</points>
<connection>
<GID>519</GID>
<name>IN_2</name></connection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-112.5,-33,-109,-33</points>
<intersection>-112.5 1</intersection>
<intersection>-109 0</intersection></hsegment></shape></wire>
<wire>
<ID>627</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106,-35.5,-106,-32</points>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-110.5,-32,-110.5,-30.5</points>
<connection>
<GID>519</GID>
<name>IN_3</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-110.5,-32,-106,-32</points>
<intersection>-110.5 1</intersection>
<intersection>-106 0</intersection></hsegment></shape></wire>
<wire>
<ID>629</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-113.5,-18.5,-113.5,-17</points>
<connection>
<GID>529</GID>
<name>OUT</name></connection>
<connection>
<GID>379</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>630</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-113.5,-24.5,-113.5,-23.5</points>
<connection>
<GID>519</GID>
<name>OUT</name></connection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-114.5,-23.5,-113.5,-23.5</points>
<intersection>-114.5 3</intersection>
<intersection>-113.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-114.5,-23.5,-114.5,-22.5</points>
<connection>
<GID>529</GID>
<name>IN_1</name></connection>
<intersection>-23.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>631</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120,-20.5,-116,-20.5</points>
<connection>
<GID>529</GID>
<name>SEL_0</name></connection>
<connection>
<GID>563</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>632</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-122,-69.5,-118,-69.5</points>
<connection>
<GID>565</GID>
<name>SEL_0</name></connection>
<connection>
<GID>566</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>661</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-97.5,-36,-93</points>
<connection>
<GID>335</GID>
<name>OUT_0</name></connection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-120,-97.5,-36,-97.5</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>-91.5 2</intersection>
<intersection>-36 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-91.5,-97.5,-91.5,-87.5</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>-97.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>662</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-111,-65,-111,-63</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>-65 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-115.5,-67.5,-115.5,-65</points>
<connection>
<GID>565</GID>
<name>OUT</name></connection>
<intersection>-65 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-115.5,-65,-111,-65</points>
<intersection>-115.5 1</intersection>
<intersection>-111 0</intersection></hsegment></shape></wire>
<wire>
<ID>668</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-111,-84.5,-103.5,-84.5</points>
<connection>
<GID>575</GID>
<name>SEL_0</name></connection>
<connection>
<GID>576</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>669</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-101,-82.5,-101,-82</points>
<connection>
<GID>575</GID>
<name>OUT</name></connection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-101,-82,-100,-82</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>-101 0</intersection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-85,-16.5,-70.5</points>
<connection>
<GID>338</GID>
<name>OUT</name></connection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32.5,-85,-16.5,-85</points>
<connection>
<GID>335</GID>
<name>IN_B_0</name></connection>
<intersection>-16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-84,-23,-70.5</points>
<connection>
<GID>339</GID>
<name>OUT</name></connection>
<intersection>-84 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-33.5,-84,-23,-84</points>
<intersection>-33.5 4</intersection>
<intersection>-23 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-33.5,-85,-33.5,-84</points>
<connection>
<GID>335</GID>
<name>IN_B_1</name></connection>
<intersection>-84 3</intersection></vsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34.5,-85,-34.5,-83</points>
<connection>
<GID>335</GID>
<name>IN_B_2</name></connection>
<intersection>-83 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-28.5,-83,-28.5,-70.5</points>
<connection>
<GID>340</GID>
<name>OUT</name></connection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-34.5,-83,-28.5,-83</points>
<intersection>-34.5 0</intersection>
<intersection>-28.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-85,-35.5,-70.5</points>
<connection>
<GID>335</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>341</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-103,-79,-102,-79</points>
<connection>
<GID>336</GID>
<name>set</name></connection>
<connection>
<GID>337</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-94,-79,-89,-79</points>
<connection>
<GID>336</GID>
<name>clear</name></connection>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>-97,-82.5,-97,-82</points>
<connection>
<GID>336</GID>
<name>clock</name></connection>
<connection>
<GID>348</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93.5,-87.5,-93.5,-74.5</points>
<intersection>-87.5 8</intersection>
<intersection>-74.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-101,-74.5,-93.5,-74.5</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>-100 11</intersection>
<intersection>-93.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-100,-87.5,-93.5,-87.5</points>
<intersection>-100 12</intersection>
<intersection>-93.5 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-100,-76,-100,-72.5</points>
<connection>
<GID>336</GID>
<name>OUT_0</name></connection>
<connection>
<GID>349</GID>
<name>N_in2</name></connection>
<intersection>-74.5 6</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>-100,-87.5,-100,-86.5</points>
<connection>
<GID>575</GID>
<name>IN_0</name></connection>
<intersection>-87.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82.5,-78.5,-81.5,-78.5</points>
<connection>
<GID>356</GID>
<name>set</name></connection>
<connection>
<GID>357</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-73.5,-78.5,-71,-78.5</points>
<connection>
<GID>356</GID>
<name>clear</name></connection>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>-76.5,-82,-76.5,-81.5</points>
<connection>
<GID>356</GID>
<name>clock</name></connection>
<connection>
<GID>359</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68,-87,-68,-73.5</points>
<intersection>-87 14</intersection>
<intersection>-73.5 15</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-78.5,-87,-68,-87</points>
<intersection>-78.5 19</intersection>
<intersection>-68 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-79.5,-73.5,-68,-73.5</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>-79.5 18</intersection>
<intersection>-68 0</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>-79.5,-75.5,-79.5,-72</points>
<connection>
<GID>356</GID>
<name>OUT_0</name></connection>
<connection>
<GID>360</GID>
<name>N_in2</name></connection>
<intersection>-73.5 15</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>-78.5,-87,-78.5,-85.5</points>
<connection>
<GID>577</GID>
<name>IN_0</name></connection>
<intersection>-87 14</intersection></vsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-114,-60,-113,-60</points>
<connection>
<GID>364</GID>
<name>set</name></connection>
<connection>
<GID>366</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105,-60,-104,-60</points>
<connection>
<GID>364</GID>
<name>clear</name></connection>
<connection>
<GID>368</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>14</ID>
<points>-108,-63.5,-108,-63</points>
<connection>
<GID>364</GID>
<name>clock</name></connection>
<connection>
<GID>370</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>692</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-102,-88,-102,-86.5</points>
<connection>
<GID>575</GID>
<name>IN_1</name></connection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-106,-88,-45.5,-88</points>
<connection>
<GID>335</GID>
<name>carry_out</name></connection>
<connection>
<GID>350</GID>
<name>N_in1</name></connection>
<intersection>-102 0</intersection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-101.5,-71.5,-101.5,-55.5</points>
<intersection>-71.5 7</intersection>
<intersection>-55.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-112,-55.5,-101.5,-55.5</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>-111 10</intersection>
<intersection>-101.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-114.5,-71.5,-101.5,-71.5</points>
<connection>
<GID>565</GID>
<name>IN_0</name></connection>
<intersection>-101.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-111,-57,-111,-53.5</points>
<connection>
<GID>364</GID>
<name>OUT_0</name></connection>
<connection>
<GID>375</GID>
<name>N_in2</name></connection>
<intersection>-55.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-115.5,-13,-114.5,-13</points>
<connection>
<GID>381</GID>
<name>OUT_0</name></connection>
<intersection>-115.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-115.5,-14,-115.5,-13</points>
<connection>
<GID>379</GID>
<name>set</name></connection>
<intersection>-13 1</intersection></vsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-107.5,-13,-104.5,-13</points>
<connection>
<GID>383</GID>
<name>OUT_0</name></connection>
<intersection>-107.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-107.5,-14,-107.5,-13</points>
<connection>
<GID>379</GID>
<name>clear</name></connection>
<intersection>-13 1</intersection></vsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59.5,-65.5,-59.5,-61.5</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<connection>
<GID>354</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53,-65.5,-53,-63.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<connection>
<GID>353</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48,-65.5,-48,-63</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<connection>
<GID>352</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-41.5,-65.5,-41.5,-64</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<connection>
<GID>351</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>12</ID>
<points>-109,-18.5,-109,-17</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<intersection>-17 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-110.5,-17,-109,-17</points>
<connection>
<GID>379</GID>
<name>clock</name></connection>
<intersection>-109 12</intersection></hsegment></shape></wire>
<wire>
<ID>702</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>-82,-83.5,-82,-69.5</points>
<connection>
<GID>577</GID>
<name>SEL_0</name></connection>
<intersection>-69.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-87.5,-69.5,-82,-69.5</points>
<connection>
<GID>578</GID>
<name>IN_0</name></connection>
<intersection>-82 4</intersection></hsegment></shape></wire>
<wire>
<ID>703</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-79.5,-81.5,-79.5,-81.5</points>
<connection>
<GID>577</GID>
<name>OUT</name></connection>
<connection>
<GID>356</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>704</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80.5,-90,-80.5,-85.5</points>
<connection>
<GID>577</GID>
<name>IN_1</name></connection>
<intersection>-90 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-102.5,-90,-45.5,-90</points>
<connection>
<GID>335</GID>
<name>overflow</name></connection>
<connection>
<GID>347</GID>
<name>N_in1</name></connection>
<intersection>-80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100.5,-24,-100.5,-8.5</points>
<intersection>-24 7</intersection>
<intersection>-8.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-115,-8.5,-100.5,-8.5</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>-113.5 11</intersection>
<intersection>-100.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-112.5,-24,-100.5,-24</points>
<intersection>-112.5 10</intersection>
<intersection>-100.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-112.5,-24,-112.5,-22.5</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<intersection>-24 7</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-113.5,-11,-113.5,-6.5</points>
<connection>
<GID>389</GID>
<name>N_in2</name></connection>
<connection>
<GID>379</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17.5,-64.5,-17.5,-45.5</points>
<connection>
<GID>338</GID>
<name>IN_1</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,-45.5,-17,-45.5</points>
<connection>
<GID>593</GID>
<name>IN_0</name></connection>
<connection>
<GID>369</GID>
<name>OUT_0</name></connection>
<intersection>-17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24,-64.5,-24,-44.5</points>
<connection>
<GID>339</GID>
<name>IN_1</name></connection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,-44.5,-17,-44.5</points>
<connection>
<GID>593</GID>
<name>IN_1</name></connection>
<connection>
<GID>369</GID>
<name>OUT_1</name></connection>
<intersection>-24 0</intersection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-64.5,-29.5,-43.5</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,-43.5,-17,-43.5</points>
<connection>
<GID>593</GID>
<name>IN_2</name></connection>
<connection>
<GID>369</GID>
<name>OUT_2</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-64.5,-36.5,-42.5</points>
<connection>
<GID>341</GID>
<name>IN_1</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,-42.5,-17,-42.5</points>
<connection>
<GID>593</GID>
<name>IN_3</name></connection>
<connection>
<GID>369</GID>
<name>OUT_3</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40.5,-74,-40.5,-71.5</points>
<connection>
<GID>351</GID>
<name>OUT</name></connection>
<connection>
<GID>371</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39.5,-85,-39.5,-80</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<connection>
<GID>371</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-47,-74.5,-47,-71.5</points>
<connection>
<GID>352</GID>
<name>OUT</name></connection>
<connection>
<GID>372</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40.5,-85,-40.5,-81.5</points>
<connection>
<GID>335</GID>
<name>IN_1</name></connection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-46,-81.5,-40.5,-81.5</points>
<intersection>-46 3</intersection>
<intersection>-40.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-46,-81.5,-46,-80.5</points>
<connection>
<GID>372</GID>
<name>OUT</name></connection>
<intersection>-81.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-41.5,-85,-41.5,-82.5</points>
<connection>
<GID>335</GID>
<name>IN_2</name></connection>
<intersection>-82.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-51,-82.5,-51,-80.5</points>
<connection>
<GID>373</GID>
<name>OUT</name></connection>
<intersection>-82.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-51,-82.5,-41.5,-82.5</points>
<intersection>-51 1</intersection>
<intersection>-41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-85,-42.5,-83.5</points>
<connection>
<GID>335</GID>
<name>IN_3</name></connection>
<intersection>-83.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-57.5,-83.5,-57.5,-80.5</points>
<connection>
<GID>374</GID>
<name>OUT</name></connection>
<intersection>-83.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,-83.5,-42.5,-83.5</points>
<intersection>-57.5 1</intersection>
<intersection>-42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-74.5,-52,-71.5</points>
<connection>
<GID>353</GID>
<name>OUT</name></connection>
<connection>
<GID>373</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58.5,-74.5,-58.5,-71.5</points>
<connection>
<GID>354</GID>
<name>OUT</name></connection>
<connection>
<GID>374</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56.5,-74.5,-56.5,-73</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60,-73,-38.5,-73</points>
<connection>
<GID>376</GID>
<name>OUT_0</name></connection>
<intersection>-56.5 0</intersection>
<intersection>-50 3</intersection>
<intersection>-45 5</intersection>
<intersection>-38.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-50,-74.5,-50,-73</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>-73 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-45,-74.5,-45,-73</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>-73 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-38.5,-74,-38.5,-73</points>
<connection>
<GID>371</GID>
<name>IN_0</name></connection>
<intersection>-73 1</intersection></vsegment></shape></wire>
<wire>
<ID>719</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-6.5,-16,-0.5</points>
<connection>
<GID>660</GID>
<name>OUT_0</name></connection>
<connection>
<GID>479</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57.5,-65.5,-57.5,-52.5</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57.5,-52.5,-10,-52.5</points>
<connection>
<GID>606</GID>
<name>IN_0</name></connection>
<intersection>-57.5 0</intersection>
<intersection>-51 7</intersection>
<intersection>-46 6</intersection>
<intersection>-39.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-39.5,-65.5,-39.5,-52.5</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-46,-65.5,-46,-52.5</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-51,-65.5,-51,-52.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34.5,-64.5,-34.5,-53.5</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-53.5,-15.5,-53.5</points>
<intersection>-34.5 0</intersection>
<intersection>-27.5 3</intersection>
<intersection>-22 7</intersection>
<intersection>-15.5 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-27.5,-64.5,-27.5,-53.5</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-15.5,-64.5,-15.5,-53.5</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>-56.5 10</intersection>
<intersection>-53.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-22,-64.5,-22,-53.5</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-15.5,-56.5,-8,-56.5</points>
<connection>
<GID>605</GID>
<name>IN_0</name></connection>
<intersection>-15.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-96,-37,-93</points>
<connection>
<GID>335</GID>
<name>OUT_1</name></connection>
<intersection>-96 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-125.5,-96,-37,-96</points>
<connection>
<GID>391</GID>
<name>IN_0</name></connection>
<intersection>-89.5 13</intersection>
<intersection>-37 0</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-89.5,-96,-89.5,-87.5</points>
<connection>
<GID>397</GID>
<name>IN_1</name></connection>
<intersection>-96 8</intersection></vsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38,-94.5,-38,-93</points>
<connection>
<GID>335</GID>
<name>OUT_2</name></connection>
<intersection>-94.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-119,-94.5,-38,-94.5</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>-87.5 13</intersection>
<intersection>-38 0</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-87.5,-94.5,-87.5,-87.5</points>
<connection>
<GID>397</GID>
<name>IN_2</name></connection>
<intersection>-94.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<hsegment>
<ID>10</ID>
<points>-125,-93,-39,-93</points>
<connection>
<GID>335</GID>
<name>OUT_3</name></connection>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<intersection>-116.5 16</intersection>
<intersection>-85.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-85.5,-93,-85.5,-87.5</points>
<connection>
<GID>397</GID>
<name>IN_3</name></connection>
<intersection>-93 10</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-116.5,-93,-116.5,-71.5</points>
<connection>
<GID>565</GID>
<name>IN_1</name></connection>
<intersection>-93 10</intersection></vsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-52,-42.5,-47,-42.5</points>
<connection>
<GID>395</GID>
<name>OUT_3</name></connection>
<connection>
<GID>369</GID>
<name>IN_3</name></connection>
<intersection>-52 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-52,-42.5,-52,-36.5</points>
<connection>
<GID>396</GID>
<name>OUT_0</name></connection>
<intersection>-42.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-52,-43.5,-47,-43.5</points>
<connection>
<GID>395</GID>
<name>OUT_2</name></connection>
<connection>
<GID>369</GID>
<name>IN_2</name></connection>
<intersection>-51 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-51,-43.5,-51,-36.5</points>
<connection>
<GID>396</GID>
<name>OUT_1</name></connection>
<intersection>-43.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-52,-44.5,-47,-44.5</points>
<connection>
<GID>395</GID>
<name>OUT_1</name></connection>
<connection>
<GID>369</GID>
<name>IN_1</name></connection>
<intersection>-50 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-50,-44.5,-50,-36.5</points>
<connection>
<GID>396</GID>
<name>OUT_2</name></connection>
<intersection>-44.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-52,-45.5,-47,-45.5</points>
<connection>
<GID>395</GID>
<name>OUT_0</name></connection>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<intersection>-49 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-49,-45.5,-49,-36.5</points>
<connection>
<GID>396</GID>
<name>OUT_3</name></connection>
<intersection>-45.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59,-42.5,-56,-42.5</points>
<connection>
<GID>395</GID>
<name>IN_3</name></connection>
<connection>
<GID>398</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-63.5,-43.5,-56,-43.5</points>
<connection>
<GID>395</GID>
<name>IN_2</name></connection>
<connection>
<GID>399</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69,-44.5,-56,-44.5</points>
<connection>
<GID>395</GID>
<name>IN_1</name></connection>
<connection>
<GID>400</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-75,-45.5,-56,-45.5</points>
<connection>
<GID>395</GID>
<name>IN_0</name></connection>
<connection>
<GID>401</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,-32.5,-49,-31</points>
<connection>
<GID>396</GID>
<name>IN_3</name></connection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-2,-45.5,-2,-25.5</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<intersection>-45.5 4</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-49,-31,-2,-31</points>
<intersection>-49 0</intersection>
<intersection>-2 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-13,-45.5,-2,-45.5</points>
<connection>
<GID>593</GID>
<name>OUT_0</name></connection>
<intersection>-2 1</intersection></hsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-44.5,-6,-25</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<intersection>-44.5 6</intersection>
<intersection>-29.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-50,-29.5,-6,-29.5</points>
<intersection>-50 4</intersection>
<intersection>-6 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-50,-32.5,-50,-29.5</points>
<connection>
<GID>396</GID>
<name>IN_2</name></connection>
<intersection>-29.5 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-13,-44.5,-6,-44.5</points>
<connection>
<GID>593</GID>
<name>OUT_1</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51,-32.5,-51,-28.5</points>
<connection>
<GID>396</GID>
<name>IN_1</name></connection>
<intersection>-28.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-51,-28.5,-10,-28.5</points>
<intersection>-51 0</intersection>
<intersection>-10 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-10,-43.5,-10,-24.5</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<intersection>-43.5 7</intersection>
<intersection>-28.5 3</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-13,-43.5,-10,-43.5</points>
<connection>
<GID>593</GID>
<name>OUT_2</name></connection>
<intersection>-10 5</intersection></hsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-32.5,-52,-26.5</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>-26.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-13,-42.5,-13,-24.5</points>
<connection>
<GID>593</GID>
<name>OUT_3</name></connection>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-52,-26.5,-13,-26.5</points>
<intersection>-52 0</intersection>
<intersection>-13 1</intersection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-50,-44,-48.5</points>
<connection>
<GID>369</GID>
<name>clock</name></connection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47.5,-50,-44,-50</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42,-48.5,-42,-48.5</points>
<connection>
<GID>407</GID>
<name>OUT_0</name></connection>
<connection>
<GID>369</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-39.5,-43,-37.5</points>
<connection>
<GID>408</GID>
<name>OUT_0</name></connection>
<connection>
<GID>369</GID>
<name>count_enable</name></connection>
<intersection>-39.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-43,-39.5,-42,-39.5</points>
<connection>
<GID>369</GID>
<name>count_up</name></connection>
<intersection>-43 0</intersection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-85.5,139,-71</points>
<connection>
<GID>432</GID>
<name>OUT</name></connection>
<intersection>-85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-85.5,139,-85.5</points>
<connection>
<GID>431</GID>
<name>IN_B_0</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,-84.5,132.5,-71</points>
<connection>
<GID>433</GID>
<name>OUT</name></connection>
<intersection>-84.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-84.5,132.5,-84.5</points>
<intersection>122 4</intersection>
<intersection>132.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>122,-85.5,122,-84.5</points>
<connection>
<GID>431</GID>
<name>IN_B_1</name></connection>
<intersection>-84.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-85.5,121,-83.5</points>
<connection>
<GID>431</GID>
<name>IN_B_2</name></connection>
<intersection>-83.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>127,-83.5,127,-71</points>
<connection>
<GID>434</GID>
<name>OUT</name></connection>
<intersection>-83.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>121,-83.5,127,-83.5</points>
<intersection>121 0</intersection>
<intersection>127 1</intersection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-85.5,120,-71</points>
<connection>
<GID>431</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>435</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47.5,-34.5,-41,-34.5</points>
<connection>
<GID>396</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>382</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-35,108,-35</points>
<connection>
<GID>419</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>384</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-66,96,-62</points>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<connection>
<GID>443</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-66,102.5,-62</points>
<connection>
<GID>438</GID>
<name>IN_0</name></connection>
<connection>
<GID>442</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-66,107.5,-62.5</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<connection>
<GID>441</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-66,114,-63</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<connection>
<GID>440</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-65,138,-46</points>
<connection>
<GID>432</GID>
<name>IN_1</name></connection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-46,139.5,-46</points>
<connection>
<GID>450</GID>
<name>OUT_0</name></connection>
<connection>
<GID>591</GID>
<name>IN_0</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-65,131.5,-45</points>
<connection>
<GID>433</GID>
<name>IN_1</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-45,139.5,-45</points>
<connection>
<GID>450</GID>
<name>OUT_1</name></connection>
<connection>
<GID>591</GID>
<name>IN_1</name></connection>
<intersection>131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-65,126,-44</points>
<connection>
<GID>434</GID>
<name>IN_1</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-44,139.5,-44</points>
<connection>
<GID>450</GID>
<name>OUT_2</name></connection>
<connection>
<GID>591</GID>
<name>IN_2</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-65,119,-43</points>
<connection>
<GID>435</GID>
<name>IN_1</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-43,139.5,-43</points>
<connection>
<GID>450</GID>
<name>OUT_3</name></connection>
<connection>
<GID>591</GID>
<name>IN_3</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-74.5,115,-72</points>
<connection>
<GID>440</GID>
<name>OUT</name></connection>
<connection>
<GID>451</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-85.5,116,-80.5</points>
<connection>
<GID>431</GID>
<name>IN_0</name></connection>
<connection>
<GID>451</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-75,108.5,-72</points>
<connection>
<GID>441</GID>
<name>OUT</name></connection>
<connection>
<GID>452</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-85.5,115,-82</points>
<connection>
<GID>431</GID>
<name>IN_1</name></connection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>109.5,-82,115,-82</points>
<intersection>109.5 4</intersection>
<intersection>115 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>109.5,-82,109.5,-81</points>
<connection>
<GID>452</GID>
<name>OUT</name></connection>
<intersection>-82 2</intersection></vsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-85.5,114,-83</points>
<connection>
<GID>431</GID>
<name>IN_2</name></connection>
<intersection>-83 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>104.5,-83,104.5,-81</points>
<connection>
<GID>453</GID>
<name>OUT</name></connection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-83,114,-83</points>
<intersection>104.5 1</intersection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-85.5,113,-84</points>
<connection>
<GID>431</GID>
<name>IN_3</name></connection>
<intersection>-84 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>98,-84,98,-81</points>
<connection>
<GID>454</GID>
<name>OUT</name></connection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>98,-84,113,-84</points>
<intersection>98 1</intersection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-75,103.5,-72</points>
<connection>
<GID>442</GID>
<name>OUT</name></connection>
<connection>
<GID>453</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>386</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-75,97,-72</points>
<connection>
<GID>443</GID>
<name>OUT</name></connection>
<connection>
<GID>454</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-75,99,-73.5</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-73.5,117,-73.5</points>
<connection>
<GID>455</GID>
<name>OUT_0</name></connection>
<intersection>99 0</intersection>
<intersection>105.5 3</intersection>
<intersection>110.5 5</intersection>
<intersection>117 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>105.5,-75,105.5,-73.5</points>
<connection>
<GID>453</GID>
<name>IN_0</name></connection>
<intersection>-73.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>110.5,-75,110.5,-73.5</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<intersection>-73.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>117,-74.5,117,-73.5</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<intersection>-73.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-66,98,-55</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98,-55,116,-55</points>
<intersection>98 0</intersection>
<intersection>104.5 7</intersection>
<intersection>109.5 6</intersection>
<intersection>116 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>116,-66,116,-55</points>
<connection>
<GID>440</GID>
<name>IN_0</name></connection>
<intersection>-56 10</intersection>
<intersection>-55 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>109.5,-66,109.5,-55</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<intersection>-55 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>104.5,-66,104.5,-55</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>116,-56,144,-56</points>
<connection>
<GID>602</GID>
<name>IN_0</name></connection>
<intersection>116 5</intersection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>-228.763,85.2289,193.165,-130.481</PageViewport>
<gate>
<ID>3</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>-123,-4.5</position>
<input>
<ID>ENABLE_0</ID>179 </input>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>84 </input>
<input>
<ID>IN_2</ID>83 </input>
<input>
<ID>IN_3</ID>82 </input>
<input>
<ID>IN_4</ID>81 </input>
<input>
<ID>IN_5</ID>80 </input>
<input>
<ID>IN_6</ID>79 </input>
<input>
<ID>IN_7</ID>78 </input>
<output>
<ID>OUT_0</ID>178 </output>
<output>
<ID>OUT_1</ID>177 </output>
<output>
<ID>OUT_2</ID>176 </output>
<output>
<ID>OUT_3</ID>130 </output>
<output>
<ID>OUT_4</ID>93 </output>
<output>
<ID>OUT_5</ID>92 </output>
<output>
<ID>OUT_6</ID>91 </output>
<output>
<ID>OUT_7</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>7</ID>
<type>DE_TO</type>
<position>-118.5,9</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I11</lparam></gate>
<gate>
<ID>9</ID>
<type>DE_TO</type>
<position>-118.5,7</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I10</lparam></gate>
<gate>
<ID>11</ID>
<type>DE_TO</type>
<position>-118.5,4.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I9</lparam></gate>
<gate>
<ID>13</ID>
<type>DE_TO</type>
<position>-118.5,2.5</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I8</lparam></gate>
<gate>
<ID>15</ID>
<type>DE_TO</type>
<position>-107.5,-1</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I7</lparam></gate>
<gate>
<ID>17</ID>
<type>DE_TO</type>
<position>-107.5,-3</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I6</lparam></gate>
<gate>
<ID>19</ID>
<type>DE_TO</type>
<position>-107.5,-5.5</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I5</lparam></gate>
<gate>
<ID>21</ID>
<type>DE_TO</type>
<position>-107.5,-7.5</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I4</lparam></gate>
<gate>
<ID>23</ID>
<type>DE_TO</type>
<position>-113.5,-10</position>
<input>
<ID>IN_0</ID>130 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I3</lparam></gate>
<gate>
<ID>25</ID>
<type>DE_TO</type>
<position>-113.5,-12</position>
<input>
<ID>IN_0</ID>176 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I2</lparam></gate>
<gate>
<ID>803</ID>
<type>DA_FROM</type>
<position>-135,-0.5</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>804</ID>
<type>DA_FROM</type>
<position>-134.5,-3</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>805</ID>
<type>DA_FROM</type>
<position>-135.5,-6</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>806</ID>
<type>DA_FROM</type>
<position>-134.5,-9</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>807</ID>
<type>DA_FROM</type>
<position>-134.5,-11</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>808</ID>
<type>DA_FROM</type>
<position>-134.5,-14</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>809</ID>
<type>DA_FROM</type>
<position>-135,-17</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>810</ID>
<type>DA_FROM</type>
<position>-135,-21</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>38</ID>
<type>DE_TO</type>
<position>-113.5,-14.5</position>
<input>
<ID>IN_0</ID>177 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I1</lparam></gate>
<gate>
<ID>812</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>-127,7.5</position>
<input>
<ID>ENABLE_0</ID>179 </input>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>45 </input>
<input>
<ID>IN_2</ID>4 </input>
<input>
<ID>IN_3</ID>701 </input>
<output>
<ID>OUT_0</ID>89 </output>
<output>
<ID>OUT_1</ID>88 </output>
<output>
<ID>OUT_2</ID>87 </output>
<output>
<ID>OUT_3</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>-113.5,-16.5</position>
<input>
<ID>IN_0</ID>178 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC I0</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>-139.5,21</position>
<input>
<ID>IN_0</ID>179 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BUS-PC</lparam></gate>
<gate>
<ID>60</ID>
<type>DA_FROM</type>
<position>-15.5,-10.5</position>
<input>
<ID>IN_0</ID>180 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I8</lparam></gate>
<gate>
<ID>61</ID>
<type>DA_FROM</type>
<position>-18,-10.5</position>
<input>
<ID>IN_0</ID>181 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I9</lparam></gate>
<gate>
<ID>62</ID>
<type>DA_FROM</type>
<position>-20.5,-10.5</position>
<input>
<ID>IN_0</ID>182 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I10</lparam></gate>
<gate>
<ID>65</ID>
<type>DA_FROM</type>
<position>-23,-10.5</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I11</lparam></gate>
<gate>
<ID>67</ID>
<type>DA_FROM</type>
<position>5,-11</position>
<input>
<ID>IN_0</ID>188 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I4</lparam></gate>
<gate>
<ID>69</ID>
<type>DA_FROM</type>
<position>2.5,-11</position>
<input>
<ID>IN_0</ID>187 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I5</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>0,-11</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I6</lparam></gate>
<gate>
<ID>74</ID>
<type>DA_FROM</type>
<position>-2.5,-11</position>
<input>
<ID>IN_0</ID>184 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I7</lparam></gate>
<gate>
<ID>275</ID>
<type>AA_TOGGLE</type>
<position>-29.5,-63</position>
<output>
<ID>OUT_0</ID>249 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>276</ID>
<type>DE_TO</type>
<position>-16.5,-63</position>
<input>
<ID>IN_0</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ck3</lparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>25.5,-10.5</position>
<input>
<ID>IN_0</ID>192 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I0</lparam></gate>
<gate>
<ID>91</ID>
<type>DA_FROM</type>
<position>23,-10.5</position>
<input>
<ID>IN_0</ID>191 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I1</lparam></gate>
<gate>
<ID>675</ID>
<type>AA_LABEL</type>
<position>20.5,109</position>
<gparam>LABEL_TEXT Program Counter</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>677</ID>
<type>AI_REGISTER12</type>
<position>54.5,-39.5</position>
<input>
<ID>IN_0</ID>649 </input>
<input>
<ID>IN_1</ID>650 </input>
<input>
<ID>IN_10</ID>659 </input>
<input>
<ID>IN_11</ID>660 </input>
<input>
<ID>IN_2</ID>651 </input>
<input>
<ID>IN_3</ID>652 </input>
<input>
<ID>IN_4</ID>653 </input>
<input>
<ID>IN_5</ID>654 </input>
<input>
<ID>IN_6</ID>655 </input>
<input>
<ID>IN_7</ID>656 </input>
<input>
<ID>IN_8</ID>657 </input>
<input>
<ID>IN_9</ID>658 </input>
<output>
<ID>OUT_0</ID>603 </output>
<output>
<ID>OUT_1</ID>602 </output>
<output>
<ID>OUT_10</ID>596 </output>
<output>
<ID>OUT_11</ID>595 </output>
<output>
<ID>OUT_2</ID>601 </output>
<output>
<ID>OUT_3</ID>604 </output>
<output>
<ID>OUT_4</ID>600 </output>
<output>
<ID>OUT_5</ID>597 </output>
<output>
<ID>OUT_6</ID>594 </output>
<output>
<ID>OUT_7</ID>599 </output>
<output>
<ID>OUT_8</ID>598 </output>
<output>
<ID>OUT_9</ID>593 </output>
<input>
<ID>clear</ID>589 </input>
<input>
<ID>clock</ID>588 </input>
<input>
<ID>count_enable</ID>592 </input>
<input>
<ID>count_up</ID>590 </input>
<input>
<ID>load</ID>591 </input>
<gparam>VALUE_BOX -2.4,-0.8,2.4,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 12</lparam>
<lparam>MAX_COUNT 4095</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>679</ID>
<type>DA_FROM</type>
<position>53.5,-51</position>
<input>
<ID>IN_0</ID>588 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Ck</lparam></gate>
<gate>
<ID>681</ID>
<type>DA_FROM</type>
<position>55.5,-53.5</position>
<input>
<ID>IN_0</ID>589 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>683</ID>
<type>EE_VDD</type>
<position>55.5,-28.5</position>
<output>
<ID>OUT_0</ID>590 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>685</ID>
<type>DA_FROM</type>
<position>48,-30</position>
<input>
<ID>IN_0</ID>591 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load PC</lparam></gate>
<gate>
<ID>687</ID>
<type>DA_FROM</type>
<position>47.5,-24.5</position>
<input>
<ID>IN_0</ID>592 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Fetch</lparam></gate>
<gate>
<ID>109</ID>
<type>DA_FROM</type>
<position>20.5,-10.5</position>
<input>
<ID>IN_0</ID>190 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I2</lparam></gate>
<gate>
<ID>689</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>103,-37.5</position>
<input>
<ID>ENABLE_0</ID>605 </input>
<input>
<ID>IN_0</ID>600 </input>
<input>
<ID>IN_1</ID>597 </input>
<input>
<ID>IN_2</ID>594 </input>
<input>
<ID>IN_3</ID>599 </input>
<input>
<ID>IN_4</ID>598 </input>
<input>
<ID>IN_5</ID>593 </input>
<input>
<ID>IN_6</ID>596 </input>
<input>
<ID>IN_7</ID>595 </input>
<output>
<ID>OUT_0</ID>634 </output>
<output>
<ID>OUT_1</ID>635 </output>
<output>
<ID>OUT_2</ID>636 </output>
<output>
<ID>OUT_3</ID>637 </output>
<output>
<ID>OUT_4</ID>638 </output>
<output>
<ID>OUT_5</ID>639 </output>
<output>
<ID>OUT_6</ID>640 </output>
<output>
<ID>OUT_7</ID>641 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>111</ID>
<type>DA_FROM</type>
<position>18,-10.5</position>
<input>
<ID>IN_0</ID>189 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PC I3</lparam></gate>
<gate>
<ID>691</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>103,-44.5</position>
<input>
<ID>ENABLE_0</ID>605 </input>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>602 </input>
<input>
<ID>IN_2</ID>601 </input>
<input>
<ID>IN_3</ID>604 </input>
<output>
<ID>OUT_0</ID>619 </output>
<output>
<ID>OUT_1</ID>620 </output>
<output>
<ID>OUT_2</ID>621 </output>
<output>
<ID>OUT_3</ID>633 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>693</ID>
<type>DA_FROM</type>
<position>99,-26</position>
<input>
<ID>IN_0</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-BUS</lparam></gate>
<gate>
<ID>694</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>69.5,-54</position>
<input>
<ID>ENABLE_0</ID>618 </input>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>602 </input>
<input>
<ID>IN_2</ID>601 </input>
<input>
<ID>IN_3</ID>604 </input>
<output>
<ID>OUT_0</ID>606 </output>
<output>
<ID>OUT_1</ID>607 </output>
<output>
<ID>OUT_2</ID>608 </output>
<output>
<ID>OUT_3</ID>609 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>115</ID>
<type>FF_GND</type>
<position>35,-26.5</position>
<output>
<ID>OUT_0</ID>193 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>695</ID>
<type>DE_TO</type>
<position>67,-61</position>
<input>
<ID>IN_0</ID>606 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 0</lparam></gate>
<gate>
<ID>696</ID>
<type>DE_TO</type>
<position>69,-61</position>
<input>
<ID>IN_0</ID>607 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 1</lparam></gate>
<gate>
<ID>697</ID>
<type>DE_TO</type>
<position>71,-61</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 2</lparam></gate>
<gate>
<ID>698</ID>
<type>DE_TO</type>
<position>73,-61</position>
<input>
<ID>IN_0</ID>609 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 3</lparam></gate>
<gate>
<ID>699</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>78.5,-54</position>
<input>
<ID>ENABLE_0</ID>618 </input>
<input>
<ID>IN_0</ID>600 </input>
<input>
<ID>IN_1</ID>597 </input>
<input>
<ID>IN_2</ID>594 </input>
<input>
<ID>IN_3</ID>599 </input>
<output>
<ID>OUT_0</ID>610 </output>
<output>
<ID>OUT_1</ID>611 </output>
<output>
<ID>OUT_2</ID>612 </output>
<output>
<ID>OUT_3</ID>613 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>700</ID>
<type>DE_TO</type>
<position>76,-61</position>
<input>
<ID>IN_0</ID>610 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 4</lparam></gate>
<gate>
<ID>701</ID>
<type>DE_TO</type>
<position>78,-61</position>
<input>
<ID>IN_0</ID>611 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 5</lparam></gate>
<gate>
<ID>702</ID>
<type>DE_TO</type>
<position>80,-61</position>
<input>
<ID>IN_0</ID>612 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 6</lparam></gate>
<gate>
<ID>703</ID>
<type>DE_TO</type>
<position>82,-61</position>
<input>
<ID>IN_0</ID>613 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 7</lparam></gate>
<gate>
<ID>704</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>88,-54</position>
<input>
<ID>ENABLE_0</ID>618 </input>
<input>
<ID>IN_0</ID>598 </input>
<input>
<ID>IN_1</ID>593 </input>
<input>
<ID>IN_2</ID>596 </input>
<input>
<ID>IN_3</ID>595 </input>
<output>
<ID>OUT_0</ID>614 </output>
<output>
<ID>OUT_1</ID>615 </output>
<output>
<ID>OUT_2</ID>616 </output>
<output>
<ID>OUT_3</ID>617 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>705</ID>
<type>DE_TO</type>
<position>85.5,-61</position>
<input>
<ID>IN_0</ID>614 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 8</lparam></gate>
<gate>
<ID>706</ID>
<type>DE_TO</type>
<position>87.5,-61</position>
<input>
<ID>IN_0</ID>615 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 9</lparam></gate>
<gate>
<ID>707</ID>
<type>DE_TO</type>
<position>89.5,-61</position>
<input>
<ID>IN_0</ID>616 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 10</lparam></gate>
<gate>
<ID>708</ID>
<type>DE_TO</type>
<position>91.5,-61</position>
<input>
<ID>IN_0</ID>617 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Addr 11</lparam></gate>
<gate>
<ID>709</ID>
<type>DA_FROM</type>
<position>94,-54</position>
<input>
<ID>IN_0</ID>618 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID PC-ADDR</lparam></gate>
<gate>
<ID>710</ID>
<type>DE_TO</type>
<position>156,-51.5</position>
<input>
<ID>IN_0</ID>645 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 15</lparam></gate>
<gate>
<ID>711</ID>
<type>DE_TO</type>
<position>152.5,-53.5</position>
<input>
<ID>IN_0</ID>644 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 14</lparam></gate>
<gate>
<ID>712</ID>
<type>DE_TO</type>
<position>149,-54</position>
<input>
<ID>IN_0</ID>643 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 13</lparam></gate>
<gate>
<ID>713</ID>
<type>DE_TO</type>
<position>145.5,-55</position>
<input>
<ID>IN_0</ID>642 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 12</lparam></gate>
<gate>
<ID>714</ID>
<type>DE_TO</type>
<position>142.5,-55.5</position>
<input>
<ID>IN_0</ID>641 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>715</ID>
<type>DE_TO</type>
<position>139,-56.5</position>
<input>
<ID>IN_0</ID>640 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>716</ID>
<type>DE_TO</type>
<position>136,-59</position>
<input>
<ID>IN_0</ID>639 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>717</ID>
<type>DE_TO</type>
<position>132.5,-60.5</position>
<input>
<ID>IN_0</ID>638 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>718</ID>
<type>DE_TO</type>
<position>107,-65.5</position>
<input>
<ID>IN_0</ID>619 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>719</ID>
<type>DE_TO</type>
<position>111,-66.5</position>
<input>
<ID>IN_0</ID>620 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>720</ID>
<type>DE_TO</type>
<position>114.5,-66.5</position>
<input>
<ID>IN_0</ID>621 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>721</ID>
<type>DE_TO</type>
<position>116.5,-66</position>
<input>
<ID>IN_0</ID>633 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>722</ID>
<type>DE_TO</type>
<position>119,-64</position>
<input>
<ID>IN_0</ID>634 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 4</lparam></gate>
<gate>
<ID>723</ID>
<type>DE_TO</type>
<position>122,-63.5</position>
<input>
<ID>IN_0</ID>635 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 5</lparam></gate>
<gate>
<ID>724</ID>
<type>DE_TO</type>
<position>124.5,-62</position>
<input>
<ID>IN_0</ID>636 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 6</lparam></gate>
<gate>
<ID>725</ID>
<type>DE_TO</type>
<position>128,-62</position>
<input>
<ID>IN_0</ID>637 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 7</lparam></gate>
<gate>
<ID>727</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>112.5,-29</position>
<input>
<ID>ENABLE_0</ID>605 </input>
<input>
<ID>IN_0</ID>646 </input>
<input>
<ID>IN_1</ID>646 </input>
<input>
<ID>IN_2</ID>646 </input>
<input>
<ID>IN_3</ID>646 </input>
<output>
<ID>OUT_0</ID>642 </output>
<output>
<ID>OUT_1</ID>643 </output>
<output>
<ID>OUT_2</ID>644 </output>
<output>
<ID>OUT_3</ID>645 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>729</ID>
<type>FF_GND</type>
<position>109.5,-32.5</position>
<output>
<ID>OUT_0</ID>646 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>734</ID>
<type>DA_FROM</type>
<position>-135,3.5</position>
<input>
<ID>IN_0</ID>53 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Bus 8</lparam></gate>
<gate>
<ID>735</ID>
<type>DA_FROM</type>
<position>-135,6</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Bus 9</lparam></gate>
<gate>
<ID>736</ID>
<type>DA_FROM</type>
<position>-135,8.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Bus 10</lparam></gate>
<gate>
<ID>737</ID>
<type>DA_FROM</type>
<position>-135,11</position>
<input>
<ID>IN_0</ID>701 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Bus 11</lparam></gate>
<gate>
<ID>739</ID>
<type>AE_FULLADDER_4BIT</type>
<position>26,-27.5</position>
<input>
<ID>IN_0</ID>192 </input>
<input>
<ID>IN_1</ID>191 </input>
<input>
<ID>IN_2</ID>190 </input>
<input>
<ID>IN_3</ID>189 </input>
<input>
<ID>IN_B_0</ID>663 </input>
<input>
<ID>IN_B_1</ID>664 </input>
<input>
<ID>IN_B_2</ID>665 </input>
<input>
<ID>IN_B_3</ID>666 </input>
<output>
<ID>OUT_0</ID>649 </output>
<output>
<ID>OUT_1</ID>650 </output>
<output>
<ID>OUT_2</ID>651 </output>
<output>
<ID>OUT_3</ID>652 </output>
<input>
<ID>carry_in</ID>193 </input>
<output>
<ID>carry_out</ID>647 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>740</ID>
<type>AE_FULLADDER_4BIT</type>
<position>6,-27.5</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>187 </input>
<input>
<ID>IN_2</ID>186 </input>
<input>
<ID>IN_3</ID>184 </input>
<input>
<ID>IN_B_0</ID>671 </input>
<input>
<ID>IN_B_1</ID>672 </input>
<input>
<ID>IN_B_2</ID>673 </input>
<input>
<ID>IN_B_3</ID>674 </input>
<output>
<ID>OUT_0</ID>653 </output>
<output>
<ID>OUT_1</ID>654 </output>
<output>
<ID>OUT_2</ID>655 </output>
<output>
<ID>OUT_3</ID>656 </output>
<input>
<ID>carry_in</ID>647 </input>
<output>
<ID>carry_out</ID>648 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>741</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-15,-27.5</position>
<input>
<ID>IN_0</ID>180 </input>
<input>
<ID>IN_1</ID>181 </input>
<input>
<ID>IN_2</ID>182 </input>
<input>
<ID>IN_3</ID>183 </input>
<input>
<ID>IN_B_0</ID>676 </input>
<input>
<ID>IN_B_1</ID>677 </input>
<input>
<ID>IN_B_2</ID>678 </input>
<input>
<ID>IN_B_3</ID>679 </input>
<output>
<ID>OUT_0</ID>657 </output>
<output>
<ID>OUT_1</ID>658 </output>
<output>
<ID>OUT_2</ID>659 </output>
<output>
<ID>OUT_3</ID>660 </output>
<input>
<ID>carry_in</ID>648 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>747</ID>
<type>AA_AND2</type>
<position>51,-20</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>667 </input>
<output>
<ID>OUT</ID>663 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>748</ID>
<type>AA_AND2</type>
<position>50.5,-15</position>
<input>
<ID>IN_0</ID>602 </input>
<input>
<ID>IN_1</ID>667 </input>
<output>
<ID>OUT</ID>664 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>749</ID>
<type>AA_AND2</type>
<position>50.5,-10</position>
<input>
<ID>IN_0</ID>601 </input>
<input>
<ID>IN_1</ID>667 </input>
<output>
<ID>OUT</ID>665 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>750</ID>
<type>AA_AND2</type>
<position>50,-5</position>
<input>
<ID>IN_0</ID>604 </input>
<input>
<ID>IN_1</ID>667 </input>
<output>
<ID>OUT</ID>666 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>752</ID>
<type>DA_FROM</type>
<position>64.5,-4</position>
<input>
<ID>IN_0</ID>667 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Offset</lparam></gate>
<gate>
<ID>760</ID>
<type>AA_AND2</type>
<position>70,1.5</position>
<input>
<ID>IN_0</ID>600 </input>
<input>
<ID>IN_1</ID>670 </input>
<output>
<ID>OUT</ID>671 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>761</ID>
<type>AA_AND2</type>
<position>69.5,6.5</position>
<input>
<ID>IN_0</ID>597 </input>
<input>
<ID>IN_1</ID>670 </input>
<output>
<ID>OUT</ID>672 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>762</ID>
<type>AA_AND2</type>
<position>69.5,11.5</position>
<input>
<ID>IN_0</ID>594 </input>
<input>
<ID>IN_1</ID>670 </input>
<output>
<ID>OUT</ID>673 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>763</ID>
<type>AA_AND2</type>
<position>69,16.5</position>
<input>
<ID>IN_0</ID>599 </input>
<input>
<ID>IN_1</ID>670 </input>
<output>
<ID>OUT</ID>674 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>764</ID>
<type>DA_FROM</type>
<position>79.5,17.5</position>
<input>
<ID>IN_0</ID>670 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Offset</lparam></gate>
<gate>
<ID>765</ID>
<type>AA_AND2</type>
<position>79.5,24</position>
<input>
<ID>IN_0</ID>598 </input>
<input>
<ID>IN_1</ID>675 </input>
<output>
<ID>OUT</ID>676 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>766</ID>
<type>AA_AND2</type>
<position>79,29</position>
<input>
<ID>IN_0</ID>593 </input>
<input>
<ID>IN_1</ID>675 </input>
<output>
<ID>OUT</ID>677 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>767</ID>
<type>AA_AND2</type>
<position>79,34</position>
<input>
<ID>IN_0</ID>596 </input>
<input>
<ID>IN_1</ID>675 </input>
<output>
<ID>OUT</ID>678 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>768</ID>
<type>AA_AND2</type>
<position>78.5,39</position>
<input>
<ID>IN_0</ID>595 </input>
<input>
<ID>IN_1</ID>675 </input>
<output>
<ID>OUT</ID>679 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>769</ID>
<type>DA_FROM</type>
<position>93,40</position>
<input>
<ID>IN_0</ID>675 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Offset</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-26.5,34,-26.5</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<connection>
<GID>739</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-131,8,-131,8.5</points>
<intersection>8 1</intersection>
<intersection>8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-131,8,-129,8</points>
<connection>
<GID>812</GID>
<name>IN_2</name></connection>
<intersection>-131 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-133,8.5,-131,8.5</points>
<connection>
<GID>736</GID>
<name>IN_0</name></connection>
<intersection>-131 0</intersection></hsegment></shape></wire>
<wire>
<ID>588</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-49,53.5,-47</points>
<connection>
<GID>677</GID>
<name>clock</name></connection>
<connection>
<GID>679</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-51.5,55.5,-47</points>
<connection>
<GID>677</GID>
<name>clear</name></connection>
<connection>
<GID>681</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>590</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-32,55.5,-29.5</points>
<connection>
<GID>677</GID>
<name>count_up</name></connection>
<connection>
<GID>683</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-32,53.5,-30</points>
<connection>
<GID>677</GID>
<name>load</name></connection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-30,53.5,-30</points>
<connection>
<GID>685</GID>
<name>IN_0</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-32,54.5,-24.5</points>
<connection>
<GID>677</GID>
<name>count_enable</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-24.5,54.5,-24.5</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-36,101,-36</points>
<connection>
<GID>689</GID>
<name>IN_5</name></connection>
<connection>
<GID>677</GID>
<name>OUT_9</name></connection>
<intersection>87.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>87.5,-52,87.5,28</points>
<connection>
<GID>704</GID>
<name>IN_1</name></connection>
<intersection>-36 1</intersection>
<intersection>28 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>82,28,87.5,28</points>
<connection>
<GID>766</GID>
<name>IN_0</name></connection>
<intersection>87.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-39,101,-39</points>
<connection>
<GID>689</GID>
<name>IN_2</name></connection>
<connection>
<GID>677</GID>
<name>OUT_6</name></connection>
<intersection>79 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>79,-52,79,10.5</points>
<connection>
<GID>699</GID>
<name>IN_2</name></connection>
<intersection>-39 1</intersection>
<intersection>10.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>72.5,10.5,79,10.5</points>
<connection>
<GID>762</GID>
<name>IN_0</name></connection>
<intersection>79 3</intersection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-34,101,-34</points>
<connection>
<GID>689</GID>
<name>IN_7</name></connection>
<connection>
<GID>677</GID>
<name>OUT_11</name></connection>
<intersection>89.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>89.5,-52,89.5,38</points>
<connection>
<GID>704</GID>
<name>IN_3</name></connection>
<intersection>-34 1</intersection>
<intersection>38 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>81.5,38,89.5,38</points>
<connection>
<GID>768</GID>
<name>IN_0</name></connection>
<intersection>89.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-35,101,-35</points>
<connection>
<GID>689</GID>
<name>IN_6</name></connection>
<connection>
<GID>677</GID>
<name>OUT_10</name></connection>
<intersection>88.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>88.5,-52,88.5,33</points>
<connection>
<GID>704</GID>
<name>IN_2</name></connection>
<intersection>-35 1</intersection>
<intersection>33 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>82,33,88.5,33</points>
<connection>
<GID>767</GID>
<name>IN_0</name></connection>
<intersection>88.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-40,101,-40</points>
<connection>
<GID>689</GID>
<name>IN_1</name></connection>
<connection>
<GID>677</GID>
<name>OUT_5</name></connection>
<intersection>78 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>78,-52,78,5.5</points>
<connection>
<GID>699</GID>
<name>IN_1</name></connection>
<intersection>-40 1</intersection>
<intersection>5.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>72.5,5.5,78,5.5</points>
<connection>
<GID>761</GID>
<name>IN_0</name></connection>
<intersection>78 3</intersection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-37,101,-37</points>
<connection>
<GID>689</GID>
<name>IN_4</name></connection>
<connection>
<GID>677</GID>
<name>OUT_8</name></connection>
<intersection>86.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>86.5,-52,86.5,23</points>
<connection>
<GID>704</GID>
<name>IN_0</name></connection>
<intersection>-37 1</intersection>
<intersection>23 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>82.5,23,86.5,23</points>
<connection>
<GID>765</GID>
<name>IN_0</name></connection>
<intersection>86.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-38,101,-38</points>
<connection>
<GID>689</GID>
<name>IN_3</name></connection>
<connection>
<GID>677</GID>
<name>OUT_7</name></connection>
<intersection>80 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>80,-52,80,15.5</points>
<connection>
<GID>699</GID>
<name>IN_3</name></connection>
<intersection>-38 1</intersection>
<intersection>15.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>72,15.5,80,15.5</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<intersection>80 3</intersection></hsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-41,101,-41</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<connection>
<GID>677</GID>
<name>OUT_4</name></connection>
<intersection>77 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77,-52,77,0.5</points>
<connection>
<GID>699</GID>
<name>IN_0</name></connection>
<intersection>-41 1</intersection>
<intersection>0.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>73,0.5,77,0.5</points>
<connection>
<GID>760</GID>
<name>IN_0</name></connection>
<intersection>77 3</intersection></hsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-44,101,-44</points>
<connection>
<GID>691</GID>
<name>IN_2</name></connection>
<intersection>59.5 10</intersection>
<intersection>70 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>70,-52,70,-11</points>
<connection>
<GID>694</GID>
<name>IN_2</name></connection>
<intersection>-44 1</intersection>
<intersection>-11 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>53.5,-11,70,-11</points>
<connection>
<GID>749</GID>
<name>IN_0</name></connection>
<intersection>70 5</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>59.5,-44,59.5,-43</points>
<connection>
<GID>677</GID>
<name>OUT_2</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-45,101,-45</points>
<connection>
<GID>691</GID>
<name>IN_1</name></connection>
<intersection>59.5 14</intersection>
<intersection>69 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>69,-52,69,-16</points>
<connection>
<GID>694</GID>
<name>IN_1</name></connection>
<intersection>-45 1</intersection>
<intersection>-16 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>53.5,-16,69,-16</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<intersection>69 5</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>59.5,-45,59.5,-44</points>
<connection>
<GID>677</GID>
<name>OUT_1</name></connection>
<intersection>-45 1</intersection></vsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-46,101,-46</points>
<connection>
<GID>691</GID>
<name>IN_0</name></connection>
<intersection>59.5 12</intersection>
<intersection>68 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>68,-52,68,-21</points>
<connection>
<GID>694</GID>
<name>IN_0</name></connection>
<intersection>-46 1</intersection>
<intersection>-21 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>54,-21,68,-21</points>
<connection>
<GID>747</GID>
<name>IN_0</name></connection>
<intersection>68 5</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>59.5,-46,59.5,-45</points>
<connection>
<GID>677</GID>
<name>OUT_0</name></connection>
<intersection>-46 1</intersection></vsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-43,101,-43</points>
<connection>
<GID>691</GID>
<name>IN_3</name></connection>
<intersection>59.5 11</intersection>
<intersection>71 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>71,-52,71,-6</points>
<connection>
<GID>694</GID>
<name>IN_3</name></connection>
<intersection>-43 1</intersection>
<intersection>-6 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>53,-6,71,-6</points>
<connection>
<GID>750</GID>
<name>IN_0</name></connection>
<intersection>71 5</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>59.5,-43,59.5,-42</points>
<connection>
<GID>677</GID>
<name>OUT_3</name></connection>
<intersection>-43 1</intersection></vsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-41.5,103,-26</points>
<connection>
<GID>689</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>691</GID>
<name>ENABLE_0</name></connection>
<intersection>-26 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>101,-26,112.5,-26</points>
<connection>
<GID>727</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>693</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-59,67,-56</points>
<connection>
<GID>695</GID>
<name>IN_0</name></connection>
<intersection>-56 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>67,-56,68,-56</points>
<connection>
<GID>694</GID>
<name>OUT_0</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-59,69,-56</points>
<connection>
<GID>696</GID>
<name>IN_0</name></connection>
<connection>
<GID>694</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-59,71,-56</points>
<connection>
<GID>697</GID>
<name>IN_0</name></connection>
<intersection>-56 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-56,71,-56</points>
<connection>
<GID>694</GID>
<name>OUT_2</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-56.5,71,-56</points>
<connection>
<GID>694</GID>
<name>OUT_3</name></connection>
<intersection>-56.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>73,-59,73,-56.5</points>
<connection>
<GID>698</GID>
<name>IN_0</name></connection>
<intersection>-56.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>71,-56.5,73,-56.5</points>
<intersection>71 0</intersection>
<intersection>73 1</intersection></hsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-59,76,-56</points>
<connection>
<GID>700</GID>
<name>IN_0</name></connection>
<intersection>-56 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>76,-56,77,-56</points>
<connection>
<GID>699</GID>
<name>OUT_0</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-59,78,-56</points>
<connection>
<GID>701</GID>
<name>IN_0</name></connection>
<connection>
<GID>699</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-59,80,-57.5</points>
<connection>
<GID>702</GID>
<name>IN_0</name></connection>
<intersection>-57.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>79,-57.5,80,-57.5</points>
<intersection>79 5</intersection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>79,-57.5,79,-56</points>
<connection>
<GID>699</GID>
<name>OUT_2</name></connection>
<intersection>-57.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>82,-59,82,-56</points>
<connection>
<GID>703</GID>
<name>IN_0</name></connection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>80,-56,82,-56</points>
<connection>
<GID>699</GID>
<name>OUT_3</name></connection>
<intersection>82 1</intersection></hsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-59,85.5,-56</points>
<connection>
<GID>705</GID>
<name>IN_0</name></connection>
<intersection>-56 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>85.5,-56,86.5,-56</points>
<connection>
<GID>704</GID>
<name>OUT_0</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-59,87.5,-56</points>
<connection>
<GID>706</GID>
<name>IN_0</name></connection>
<connection>
<GID>704</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-59,89.5,-56</points>
<connection>
<GID>707</GID>
<name>IN_0</name></connection>
<intersection>-56 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>88.5,-56,89.5,-56</points>
<connection>
<GID>704</GID>
<name>OUT_2</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-56.5,89.5,-56</points>
<connection>
<GID>704</GID>
<name>OUT_3</name></connection>
<intersection>-56.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>91.5,-59,91.5,-56.5</points>
<connection>
<GID>708</GID>
<name>IN_0</name></connection>
<intersection>-56.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-56.5,91.5,-56.5</points>
<intersection>89.5 0</intersection>
<intersection>91.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72.5,-54,92,-54</points>
<connection>
<GID>694</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>699</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>704</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>709</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-46,107,-46</points>
<connection>
<GID>691</GID>
<name>OUT_0</name></connection>
<intersection>107 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>107,-63.5,107,-46</points>
<connection>
<GID>718</GID>
<name>IN_0</name></connection>
<intersection>-46 1</intersection></vsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-64.5,111,-45</points>
<connection>
<GID>719</GID>
<name>IN_0</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-45,111,-45</points>
<connection>
<GID>691</GID>
<name>OUT_1</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-64.5,114.5,-44</points>
<connection>
<GID>720</GID>
<name>IN_0</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-44,114.5,-44</points>
<connection>
<GID>691</GID>
<name>OUT_2</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-131,6,-131,7</points>
<intersection>6 2</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-131,7,-129,7</points>
<connection>
<GID>812</GID>
<name>IN_1</name></connection>
<intersection>-131 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-133,6,-131,6</points>
<connection>
<GID>735</GID>
<name>IN_0</name></connection>
<intersection>-131 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-130,3.5,-130,6</points>
<intersection>3.5 2</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-130,6,-129,6</points>
<connection>
<GID>812</GID>
<name>IN_0</name></connection>
<intersection>-130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-133,3.5,-130,3.5</points>
<connection>
<GID>734</GID>
<name>IN_0</name></connection>
<intersection>-130 0</intersection></hsegment></shape></wire>
<wire>
<ID>633</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-64,116.5,-43</points>
<connection>
<GID>721</GID>
<name>IN_0</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-43,116.5,-43</points>
<connection>
<GID>691</GID>
<name>OUT_3</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>634</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-62,119,-41</points>
<connection>
<GID>722</GID>
<name>IN_0</name></connection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-41,119,-41</points>
<connection>
<GID>689</GID>
<name>OUT_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>635</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-61.5,122,-40</points>
<connection>
<GID>723</GID>
<name>IN_0</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-40,122,-40</points>
<connection>
<GID>689</GID>
<name>OUT_1</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27.5,-63,-18.5,-63</points>
<connection>
<GID>275</GID>
<name>OUT_0</name></connection>
<connection>
<GID>276</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>636</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-60,124.5,-39</points>
<connection>
<GID>724</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-39,124.5,-39</points>
<connection>
<GID>689</GID>
<name>OUT_2</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>637</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-60,128,-38</points>
<connection>
<GID>725</GID>
<name>IN_0</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-38,128,-38</points>
<connection>
<GID>689</GID>
<name>OUT_3</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>638</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,-58.5,132.5,-37</points>
<connection>
<GID>717</GID>
<name>IN_0</name></connection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-37,132.5,-37</points>
<connection>
<GID>689</GID>
<name>OUT_4</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>639</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-57,136,-36</points>
<connection>
<GID>716</GID>
<name>IN_0</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-36,136,-36</points>
<connection>
<GID>689</GID>
<name>OUT_5</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-54.5,139,-35</points>
<connection>
<GID>715</GID>
<name>IN_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-35,139,-35</points>
<connection>
<GID>689</GID>
<name>OUT_6</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>641</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-53.5,142.5,-34</points>
<connection>
<GID>714</GID>
<name>IN_0</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-34,142.5,-34</points>
<connection>
<GID>689</GID>
<name>OUT_7</name></connection>
<intersection>142.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>642</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-53,145.5,-30.5</points>
<connection>
<GID>713</GID>
<name>IN_0</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-30.5,145.5,-30.5</points>
<connection>
<GID>727</GID>
<name>OUT_0</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>643</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,-52,149,-29.5</points>
<connection>
<GID>712</GID>
<name>IN_0</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-29.5,149,-29.5</points>
<connection>
<GID>727</GID>
<name>OUT_1</name></connection>
<intersection>149 0</intersection></hsegment></shape></wire>
<wire>
<ID>644</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152.5,-51.5,152.5,-28.5</points>
<connection>
<GID>711</GID>
<name>IN_0</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-28.5,152.5,-28.5</points>
<connection>
<GID>727</GID>
<name>OUT_2</name></connection>
<intersection>152.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>645</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-49.5,156,-27.5</points>
<connection>
<GID>710</GID>
<name>IN_0</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-27.5,156,-27.5</points>
<connection>
<GID>727</GID>
<name>OUT_3</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>646</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-31.5,109.5,-30.5</points>
<connection>
<GID>729</GID>
<name>OUT_0</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-30.5,110.5,-30.5</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<intersection>109.5 0</intersection>
<intersection>110.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110.5,-30.5,110.5,-27.5</points>
<connection>
<GID>727</GID>
<name>IN_3</name></connection>
<connection>
<GID>727</GID>
<name>IN_2</name></connection>
<connection>
<GID>727</GID>
<name>IN_1</name></connection>
<intersection>-30.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>647</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-26.5,18,-26.5</points>
<connection>
<GID>739</GID>
<name>carry_out</name></connection>
<connection>
<GID>740</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>648</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7,-26.5,-2,-26.5</points>
<connection>
<GID>740</GID>
<name>carry_out</name></connection>
<connection>
<GID>741</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>649</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-45,27.5,-31.5</points>
<connection>
<GID>739</GID>
<name>OUT_0</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-45,49.5,-45</points>
<connection>
<GID>677</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>650</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-44,26.5,-31.5</points>
<connection>
<GID>739</GID>
<name>OUT_1</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-44,49.5,-44</points>
<connection>
<GID>677</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>651</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-43,25.5,-31.5</points>
<connection>
<GID>739</GID>
<name>OUT_2</name></connection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-43,49.5,-43</points>
<connection>
<GID>677</GID>
<name>IN_2</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>652</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-42,24.5,-31.5</points>
<connection>
<GID>739</GID>
<name>OUT_3</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-42,49.5,-42</points>
<connection>
<GID>677</GID>
<name>IN_3</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>653</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-41,7.5,-31.5</points>
<connection>
<GID>740</GID>
<name>OUT_0</name></connection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,-41,49.5,-41</points>
<connection>
<GID>677</GID>
<name>IN_4</name></connection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>654</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-40,6.5,-31.5</points>
<connection>
<GID>740</GID>
<name>OUT_1</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-40,49.5,-40</points>
<connection>
<GID>677</GID>
<name>IN_5</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>655</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-39,5.5,-31.5</points>
<connection>
<GID>740</GID>
<name>OUT_2</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,-39,49.5,-39</points>
<connection>
<GID>677</GID>
<name>IN_6</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>656</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-38,4.5,-31.5</points>
<connection>
<GID>740</GID>
<name>OUT_3</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4.5,-38,49.5,-38</points>
<connection>
<GID>677</GID>
<name>IN_7</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>657</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-37,-13.5,-31.5</points>
<connection>
<GID>741</GID>
<name>OUT_0</name></connection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13.5,-37,49.5,-37</points>
<connection>
<GID>677</GID>
<name>IN_8</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-131,-1,-131,-0.5</points>
<intersection>-1 2</intersection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,-0.5,-131,-0.5</points>
<connection>
<GID>803</GID>
<name>IN_0</name></connection>
<intersection>-131 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-131,-1,-125,-1</points>
<connection>
<GID>3</GID>
<name>IN_7</name></connection>
<intersection>-131 0</intersection></hsegment></shape></wire>
<wire>
<ID>658</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-36,-14.5,-31.5</points>
<connection>
<GID>741</GID>
<name>OUT_1</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-36,49.5,-36</points>
<connection>
<GID>677</GID>
<name>IN_9</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-131.5,-3,-131.5,-2</points>
<intersection>-3 1</intersection>
<intersection>-2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-132.5,-3,-131.5,-3</points>
<connection>
<GID>804</GID>
<name>IN_0</name></connection>
<intersection>-131.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-131.5,-2,-125,-2</points>
<connection>
<GID>3</GID>
<name>IN_6</name></connection>
<intersection>-131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>659</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-35,-15.5,-31.5</points>
<connection>
<GID>741</GID>
<name>OUT_2</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15.5,-35,49.5,-35</points>
<connection>
<GID>677</GID>
<name>IN_10</name></connection>
<intersection>-15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-131,-6,-131,-3</points>
<intersection>-6 1</intersection>
<intersection>-3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133.5,-6,-131,-6</points>
<connection>
<GID>805</GID>
<name>IN_0</name></connection>
<intersection>-131 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-131,-3,-125,-3</points>
<connection>
<GID>3</GID>
<name>IN_5</name></connection>
<intersection>-131 0</intersection></hsegment></shape></wire>
<wire>
<ID>660</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-34,-16.5,-31.5</points>
<connection>
<GID>741</GID>
<name>OUT_3</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16.5,-34,49.5,-34</points>
<connection>
<GID>677</GID>
<name>IN_11</name></connection>
<intersection>-16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-129.5,-9,-129.5,-4</points>
<intersection>-9 1</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-132.5,-9,-129.5,-9</points>
<connection>
<GID>806</GID>
<name>IN_0</name></connection>
<intersection>-129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-129.5,-4,-125,-4</points>
<connection>
<GID>3</GID>
<name>IN_4</name></connection>
<intersection>-129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-129,-11,-129,-5</points>
<intersection>-11 1</intersection>
<intersection>-5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-132.5,-11,-129,-11</points>
<connection>
<GID>807</GID>
<name>IN_0</name></connection>
<intersection>-129 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-129,-5,-125,-5</points>
<connection>
<GID>3</GID>
<name>IN_3</name></connection>
<intersection>-129 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-128.5,-14,-128.5,-6</points>
<intersection>-14 2</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-128.5,-6,-125,-6</points>
<connection>
<GID>3</GID>
<name>IN_2</name></connection>
<intersection>-128.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-132.5,-14,-128.5,-14</points>
<connection>
<GID>808</GID>
<name>IN_0</name></connection>
<intersection>-128.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-23.5,31,-20</points>
<connection>
<GID>739</GID>
<name>IN_B_0</name></connection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-20,48,-20</points>
<connection>
<GID>747</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-127.5,-17,-127.5,-7</points>
<intersection>-17 2</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-127.5,-7,-125,-7</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>-127.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-133,-17,-127.5,-17</points>
<connection>
<GID>809</GID>
<name>IN_0</name></connection>
<intersection>-127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>664</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-23.5,30,-15</points>
<connection>
<GID>739</GID>
<name>IN_B_1</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-15,47.5,-15</points>
<connection>
<GID>748</GID>
<name>OUT</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-126.5,-21,-126.5,-8</points>
<intersection>-21 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,-21,-126.5,-21</points>
<connection>
<GID>810</GID>
<name>IN_0</name></connection>
<intersection>-126.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-126.5,-8,-125,-8</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>-126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>665</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-23.5,29,-10</points>
<connection>
<GID>739</GID>
<name>IN_B_2</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-10,47.5,-10</points>
<connection>
<GID>749</GID>
<name>OUT</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-125,9,-120.5,9</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<connection>
<GID>812</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-23.5,28,-5</points>
<connection>
<GID>739</GID>
<name>IN_B_3</name></connection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-5,47,-5</points>
<connection>
<GID>750</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-122,7,-122,8</points>
<intersection>7 2</intersection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-125,8,-122,8</points>
<connection>
<GID>812</GID>
<name>OUT_2</name></connection>
<intersection>-122 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-122,7,-120.5,7</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>-122 0</intersection></hsegment></shape></wire>
<wire>
<ID>667</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>53,-4,62.5,-4</points>
<connection>
<GID>750</GID>
<name>IN_1</name></connection>
<connection>
<GID>752</GID>
<name>IN_0</name></connection>
<intersection>54.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54.5,-19,54.5,-4</points>
<intersection>-19 8</intersection>
<intersection>-14 5</intersection>
<intersection>-9 6</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>53.5,-14,54.5,-14</points>
<connection>
<GID>748</GID>
<name>IN_1</name></connection>
<intersection>54.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>53.5,-9,54.5,-9</points>
<connection>
<GID>749</GID>
<name>IN_1</name></connection>
<intersection>54.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>54,-19,54.5,-19</points>
<connection>
<GID>747</GID>
<name>IN_1</name></connection>
<intersection>54.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-122.5,4.5,-122.5,7</points>
<intersection>4.5 2</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-125,7,-122.5,7</points>
<connection>
<GID>812</GID>
<name>OUT_1</name></connection>
<intersection>-122.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-122.5,4.5,-120.5,4.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>-122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-123,2.5,-123,6</points>
<intersection>2.5 2</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-125,6,-123,6</points>
<connection>
<GID>812</GID>
<name>OUT_0</name></connection>
<intersection>-123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-123,2.5,-120.5,2.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>-123 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-121,-1,-109.5,-1</points>
<connection>
<GID>3</GID>
<name>OUT_7</name></connection>
<connection>
<GID>15</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>670</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>72,17.5,77.5,17.5</points>
<connection>
<GID>763</GID>
<name>IN_1</name></connection>
<connection>
<GID>764</GID>
<name>IN_0</name></connection>
<intersection>73.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>73.5,2.5,73.5,17.5</points>
<intersection>2.5 8</intersection>
<intersection>7.5 5</intersection>
<intersection>12.5 6</intersection>
<intersection>17.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>72.5,7.5,73.5,7.5</points>
<connection>
<GID>761</GID>
<name>IN_1</name></connection>
<intersection>73.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>72.5,12.5,73.5,12.5</points>
<connection>
<GID>762</GID>
<name>IN_1</name></connection>
<intersection>73.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>73,2.5,73.5,2.5</points>
<connection>
<GID>760</GID>
<name>IN_1</name></connection>
<intersection>73.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110.5,-3,-110.5,-2</points>
<intersection>-3 2</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-121,-2,-110.5,-2</points>
<connection>
<GID>3</GID>
<name>OUT_6</name></connection>
<intersection>-110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-110.5,-3,-109.5,-3</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>-110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>671</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-23.5,11,1.5</points>
<connection>
<GID>740</GID>
<name>IN_B_0</name></connection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,1.5,67,1.5</points>
<connection>
<GID>760</GID>
<name>OUT</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-111.5,-5.5,-111.5,-3</points>
<intersection>-5.5 2</intersection>
<intersection>-3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-121,-3,-111.5,-3</points>
<connection>
<GID>3</GID>
<name>OUT_5</name></connection>
<intersection>-111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-111.5,-5.5,-109.5,-5.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>672</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-23.5,10,6.5</points>
<connection>
<GID>740</GID>
<name>IN_B_1</name></connection>
<intersection>6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,6.5,66.5,6.5</points>
<connection>
<GID>761</GID>
<name>OUT</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-112.5,-7.5,-112.5,-4</points>
<intersection>-7.5 1</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-112.5,-7.5,-109.5,-7.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-112.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121,-4,-112.5,-4</points>
<connection>
<GID>3</GID>
<name>OUT_4</name></connection>
<intersection>-112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>673</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-23.5,9,11.5</points>
<connection>
<GID>740</GID>
<name>IN_B_2</name></connection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,11.5,66.5,11.5</points>
<connection>
<GID>762</GID>
<name>OUT</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>674</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-23.5,8,16.5</points>
<connection>
<GID>740</GID>
<name>IN_B_3</name></connection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,16.5,66,16.5</points>
<connection>
<GID>763</GID>
<name>OUT</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>675</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>81.5,40,91,40</points>
<connection>
<GID>768</GID>
<name>IN_1</name></connection>
<connection>
<GID>769</GID>
<name>IN_0</name></connection>
<intersection>83 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>83,25,83,40</points>
<intersection>25 8</intersection>
<intersection>30 5</intersection>
<intersection>35 6</intersection>
<intersection>40 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>82,30,83,30</points>
<connection>
<GID>766</GID>
<name>IN_1</name></connection>
<intersection>83 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>82,35,83,35</points>
<connection>
<GID>767</GID>
<name>IN_1</name></connection>
<intersection>83 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>82.5,25,83,25</points>
<connection>
<GID>765</GID>
<name>IN_1</name></connection>
<intersection>83 3</intersection></hsegment></shape></wire>
<wire>
<ID>676</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-23.5,-10,24</points>
<connection>
<GID>741</GID>
<name>IN_B_0</name></connection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10,24,76.5,24</points>
<connection>
<GID>765</GID>
<name>OUT</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>677</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-23.5,-11,29</points>
<connection>
<GID>741</GID>
<name>IN_B_1</name></connection>
<intersection>29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11,29,76,29</points>
<connection>
<GID>766</GID>
<name>OUT</name></connection>
<intersection>-11 0</intersection></hsegment></shape></wire>
<wire>
<ID>678</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-23.5,-12,34</points>
<connection>
<GID>741</GID>
<name>IN_B_2</name></connection>
<intersection>34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,34,76,34</points>
<connection>
<GID>767</GID>
<name>OUT</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>679</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,-23.5,-13,39</points>
<connection>
<GID>741</GID>
<name>IN_B_3</name></connection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,39,75.5,39</points>
<connection>
<GID>768</GID>
<name>OUT</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>701</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-131,9,-131,11</points>
<intersection>9 2</intersection>
<intersection>11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-133,11,-131,11</points>
<connection>
<GID>737</GID>
<name>IN_0</name></connection>
<intersection>-131 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-131,9,-129,9</points>
<connection>
<GID>812</GID>
<name>IN_3</name></connection>
<intersection>-131 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-115.5,-10,-115.5,-5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-121,-5,-115.5,-5</points>
<connection>
<GID>3</GID>
<name>OUT_3</name></connection>
<intersection>-115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-116.5,-12,-116.5,-6</points>
<intersection>-12 1</intersection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-116.5,-12,-115.5,-12</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121,-6,-116.5,-6</points>
<connection>
<GID>3</GID>
<name>OUT_2</name></connection>
<intersection>-116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-117.5,-14.5,-117.5,-7</points>
<intersection>-14.5 1</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-117.5,-14.5,-115.5,-14.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121,-7,-117.5,-7</points>
<connection>
<GID>3</GID>
<name>OUT_1</name></connection>
<intersection>-117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-118.5,-16.5,-118.5,-8</points>
<intersection>-16.5 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-118.5,-16.5,-115.5,-16.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>-118.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121,-8,-118.5,-8</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-127,0.5,-127,21</points>
<connection>
<GID>812</GID>
<name>ENABLE_0</name></connection>
<intersection>0.5 2</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-137.5,21,-127,21</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-127 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-127,0.5,-123,0.5</points>
<connection>
<GID>3</GID>
<name>ENABLE_0</name></connection>
<intersection>-127 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,-23.5,-17,-18</points>
<connection>
<GID>741</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-15.5,-18,-15.5,-12.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-17,-18,-15.5,-18</points>
<intersection>-17 0</intersection>
<intersection>-15.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18,-23.5,-18,-12.5</points>
<connection>
<GID>741</GID>
<name>IN_1</name></connection>
<connection>
<GID>61</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19,-23.5,-19,-18</points>
<connection>
<GID>741</GID>
<name>IN_2</name></connection>
<intersection>-18 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-20.5,-18,-20.5,-12.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-20.5,-18,-19,-18</points>
<intersection>-20.5 1</intersection>
<intersection>-19 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,-23.5,-20,-19</points>
<connection>
<GID>741</GID>
<name>IN_3</name></connection>
<intersection>-19 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-23,-19,-23,-12.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-23,-19,-20,-19</points>
<intersection>-23 1</intersection>
<intersection>-20 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-23.5,1,-22</points>
<connection>
<GID>740</GID>
<name>IN_3</name></connection>
<intersection>-22 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-2.5,-22,-2.5,-13</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-2.5,-22,1,-22</points>
<intersection>-2.5 1</intersection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-23.5,2,-21</points>
<connection>
<GID>740</GID>
<name>IN_2</name></connection>
<intersection>-21 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-7.30078e-008,-21,-7.30078e-008,-13</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-7.30078e-008,-21,2,-21</points>
<intersection>-7.30078e-008 1</intersection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-23.5,3,-18</points>
<connection>
<GID>740</GID>
<name>IN_1</name></connection>
<intersection>-18 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>2.5,-18,2.5,-13</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>2.5,-18,3,-18</points>
<intersection>2.5 1</intersection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-23.5,4,-18</points>
<connection>
<GID>740</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>5,-18,5,-13</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>4,-18,5,-18</points>
<intersection>4 0</intersection>
<intersection>5 1</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-23.5,21,-20.5</points>
<connection>
<GID>739</GID>
<name>IN_3</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>18,-20.5,18,-12.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>18,-20.5,21,-20.5</points>
<intersection>18 1</intersection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-23.5,22,-18</points>
<connection>
<GID>739</GID>
<name>IN_2</name></connection>
<intersection>-18 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>20.5,-18,20.5,-12.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>20.5,-18,22,-18</points>
<intersection>20.5 1</intersection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-23.5,23,-12.5</points>
<connection>
<GID>739</GID>
<name>IN_1</name></connection>
<connection>
<GID>91</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-23.5,24,-18</points>
<connection>
<GID>739</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>25.5,-18,25.5,-12.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>24,-18,25.5,-18</points>
<intersection>24 0</intersection>
<intersection>25.5 1</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>-23.4529,1897.92,1754.55,988.92</PageViewport></page 6>
<page 7>
<PageViewport>-23.4529,1897.92,1754.55,988.92</PageViewport></page 7>
<page 8>
<PageViewport>-23.4529,1897.92,1754.55,988.92</PageViewport></page 8>
<page 9>
<PageViewport>-23.4529,1897.92,1754.55,988.92</PageViewport></page 9></circuit>