<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>3,0,84.6,-90</PageViewport>
<gate>
<ID>4</ID>
<type>DE_TO</type>
<position>12.5,-12</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input A</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>5,-12</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>DE_TO</type>
<position>13,-21</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input B</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>5,-21</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>DA_FROM</type>
<position>37,-11.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Input A</lparam></gate>
<gate>
<ID>13</ID>
<type>DA_FROM</type>
<position>37,-22.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Input B</lparam></gate>
<gate>
<ID>17</ID>
<type>BE_NOR2</type>
<position>45.5,-12.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>BE_NOR2</type>
<position>45.5,-21.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>GA_LED</type>
<position>62,-12.5</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>62,-21.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>5.5,-37</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>DE_TO</type>
<position>15.5,-37</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Data</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>5.5,-43</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>DE_TO</type>
<position>16,-43</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Enable</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>32.5,-37</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Data</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>34.5,-47</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Enable</lparam></gate>
<gate>
<ID>35</ID>
<type>AE_SMALL_INVERTER</type>
<position>41,-37</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_AND2</type>
<position>50.5,-36</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>50.5,-46</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>BE_NOR2</type>
<position>64.5,-37</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>GA_LED</type>
<position>76.5,-37</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>BE_NOR2</type>
<position>64.5,-45</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>GA_LED</type>
<position>76.5,-45</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-12,10.5,-12</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-21,11,-21</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-11.5,42.5,-11.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-22.5,42.5,-22.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-12.5,61,-12.5</points>
<connection>
<GID>21</GID>
<name>N_in0</name></connection>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>56.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>56.5,-27.5,56.5,-12.5</points>
<intersection>-27.5 5</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>42.5,-27.5,56.5,-27.5</points>
<intersection>42.5 6</intersection>
<intersection>56.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>42.5,-27.5,42.5,-20.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-27.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-21.5,61,-21.5</points>
<connection>
<GID>23</GID>
<name>N_in0</name></connection>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>54 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>54,-21.5,54,-18</points>
<intersection>-21.5 1</intersection>
<intersection>-18 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>42.5,-18,54,-18</points>
<intersection>42.5 12</intersection>
<intersection>54 10</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>42.5,-18,42.5,-13.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>-18 11</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-37,13.5,-37</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>7.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>7.5,-37,7.5,-37</points>
<intersection>-37 1</intersection>
<intersection>-37 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>7.5,-37,7.5,-37</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>7.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-43,14,-43</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-37,39,-37</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>37 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37,-45,37,-37</points>
<intersection>-45 4</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37,-45,47.5,-45</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>37 3</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-37,47.5,-37</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36.5,-47,47.5,-47</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>43.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>43.5,-47,43.5,-35</points>
<intersection>-47 1</intersection>
<intersection>-35 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>43.5,-35,47.5,-35</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>43.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-36,61.5,-36</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<connection>
<GID>37</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>67.5,-37,75.5,-37</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<connection>
<GID>41</GID>
<name>N_in0</name></connection>
<intersection>71 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>71,-41,71,-37</points>
<intersection>-41 6</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>61.5,-41,71,-41</points>
<intersection>61.5 7</intersection>
<intersection>71 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>61.5,-44,61.5,-41</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-41 6</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-46,61.5,-46</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<connection>
<GID>38</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-42,72.5,-42</points>
<intersection>57.5 3</intersection>
<intersection>72.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>57.5,-42,57.5,-38</points>
<intersection>-42 1</intersection>
<intersection>-38 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>57.5,-38,61.5,-38</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>57.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>72.5,-45,72.5,-42</points>
<intersection>-45 7</intersection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>67.5,-45,75.5,-45</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<connection>
<GID>43</GID>
<name>N_in0</name></connection>
<intersection>72.5 5</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,81.6,-90</PageViewport></page 1>
<page 2>
<PageViewport>0,0,81.6,-90</PageViewport></page 2>
<page 3>
<PageViewport>0,0,81.6,-90</PageViewport></page 3>
<page 4>
<PageViewport>0,0,81.6,-90</PageViewport></page 4>
<page 5>
<PageViewport>0,0,81.6,-90</PageViewport></page 5>
<page 6>
<PageViewport>0,0,81.6,-90</PageViewport></page 6>
<page 7>
<PageViewport>0,0,81.6,-90</PageViewport></page 7>
<page 8>
<PageViewport>0,0,81.6,-90</PageViewport></page 8>
<page 9>
<PageViewport>0,0,81.6,-90</PageViewport></page 9></circuit>