<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-81.9752,-85.0408,151.282,-342.309</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>-8.5,-74.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2</ID>
<type>DE_TO</type>
<position>1,-74.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Data2</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>-9.5,-83.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>DE_TO</type>
<position>17.5,31.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input A</lparam></gate>
<gate>
<ID>5</ID>
<type>DE_TO</type>
<position>-1,-83.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Enable2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>10,31.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>DA_FROM</type>
<position>27.5,-74</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Data2</lparam></gate>
<gate>
<ID>8</ID>
<type>DE_TO</type>
<position>18,22.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input B</lparam></gate>
<gate>
<ID>9</ID>
<type>DA_FROM</type>
<position>29.5,-84</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Enable2</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>10,22.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>11</ID>
<type>AE_SMALL_INVERTER</type>
<position>33.5,-78.5</position>
<input>
<ID>IN_0</ID>35 </input>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>DA_FROM</type>
<position>42,32</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Input A</lparam></gate>
<gate>
<ID>13</ID>
<type>DA_FROM</type>
<position>42,21</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Input B</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND2</type>
<position>45.5,-73</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_AND2</type>
<position>47.5,-83</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>BE_NOR2</type>
<position>59.5,-74</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>BE_NOR2</type>
<position>50.5,31</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>70.5,-67</position>
<input>
<ID>N_in2</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>BE_NOR2</type>
<position>50.5,22</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>BE_NOR2</type>
<position>59.5,-82</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>GA_LED</type>
<position>67,31</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>70,-87.5</position>
<input>
<ID>N_in3</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>67,22</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>80.5,-73</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>2.5,2</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_AND2</type>
<position>80.5,-82.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>DE_TO</type>
<position>12.5,2</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Data</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>2.5,-4</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>DE_TO</type>
<position>13,-4</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Enable</lparam></gate>
<gate>
<ID>30</ID>
<type>DE_TO</type>
<position>2.5,-127</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Enable3</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>29.5,2</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Data</lparam></gate>
<gate>
<ID>32</ID>
<type>DE_TO</type>
<position>1,-149.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Data3</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>31.5,-8</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Enable</lparam></gate>
<gate>
<ID>35</ID>
<type>AE_SMALL_INVERTER</type>
<position>38,2</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AE_SMALL_INVERTER</type>
<position>36,-84</position>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_AND2</type>
<position>47.5,3</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>47.5,-7</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>BE_NOR2</type>
<position>93,-73</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>BE_NOR2</type>
<position>61.5,2</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>GA_LED</type>
<position>73.5,2</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>BE_NOR2</type>
<position>61.5,-6</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>GA_LED</type>
<position>73.5,-6</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>BE_NOR2</type>
<position>93.5,-81.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>-10,-127</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>-10,-149.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>110.5,-73</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>DA_FROM</type>
<position>35.5,-137.5</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Enable3</lparam></gate>
<gate>
<ID>50</ID>
<type>DA_FROM</type>
<position>35,-127</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Data3</lparam></gate>
<gate>
<ID>52</ID>
<type>GA_LED</type>
<position>110,-81.5</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AE_SMALL_INVERTER</type>
<position>45,-137.5</position>
<input>
<ID>IN_0</ID>20 </input>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>55</ID>
<type>BA_NAND2</type>
<position>57.5,-136.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>BA_NAND2</type>
<position>57,-128</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>BA_NAND2</type>
<position>71,-128</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>55,-57</position>
<gparam>LABEL_TEXT Master-Slave circuit</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>BA_NAND2</type>
<position>71.5,-136.5</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>GA_LED</type>
<position>75.5,-121.5</position>
<input>
<ID>N_in2</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>75.5,-144</position>
<input>
<ID>N_in0</ID>29 </input>
<input>
<ID>N_in1</ID>29 </input>
<input>
<ID>N_in3</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>BA_NAND2</type>
<position>84.5,-128</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>BA_NAND2</type>
<position>85.5,-136.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>BA_NAND2</type>
<position>102,-127.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>BA_NAND2</type>
<position>102,-137</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>GA_LED</type>
<position>115.5,-127.5</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>GA_LED</type>
<position>116,-137.5</position>
<input>
<ID>N_in0</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>57.5,-109</position>
<gparam>LABEL_TEXT Master-slave Only NAND and Inverter</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>29.5,-181</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Data4</lparam></gate>
<gate>
<ID>72</ID>
<type>DA_FROM</type>
<position>29.5,-194.5</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Enable4</lparam></gate>
<gate>
<ID>73</ID>
<type>DE_TO</type>
<position>-1.5,-195</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Enable4</lparam></gate>
<gate>
<ID>74</ID>
<type>DE_TO</type>
<position>-0.5,-173.5</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Data4</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_TOGGLE</type>
<position>-16.5,-195</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_TOGGLE</type>
<position>-12.5,-173.5</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_TOGGLE</type>
<position>-16,-207.5</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>82</ID>
<type>DE_TO</type>
<position>2,-207.5</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>84</ID>
<type>DA_FROM</type>
<position>29,-187</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_AND3</type>
<position>54.5,-180.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>66 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_AND3</type>
<position>54.5,-194.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>66 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>88</ID>
<type>BE_NOR2</type>
<position>69.5,-181.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>BE_NOR2</type>
<position>69.5,-193.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>90</ID>
<type>AE_SMALL_INVERTER</type>
<position>40,-181</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>angle 0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>92</ID>
<type>GA_LED</type>
<position>77.5,-171</position>
<input>
<ID>N_in2</ID>57 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>GA_LED</type>
<position>77.5,-200.5</position>
<input>
<ID>N_in3</ID>58 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_AND2</type>
<position>98,-182</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_AND2</type>
<position>98.5,-194.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>100</ID>
<type>BE_NOR2</type>
<position>119.5,-182</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>BE_NOR2</type>
<position>121,-195</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>GA_LED</type>
<position>151,-182</position>
<input>
<ID>N_in3</ID>61 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>GA_LED</type>
<position>151.5,-195</position>
<input>
<ID>N_in0</ID>62 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AE_SMALL_INVERTER</type>
<position>42,-187</position>
<input>
<ID>IN_0</ID>65 </input>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>62.5,-157.5</position>
<gparam>LABEL_TEXT Master-slave with clock</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,31.5,15.5,31.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,22.5,16,22.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-74.5,-1,-74.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-6.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-6.5,-74.5,-6.5,-74.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>-74.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,32,47.5,32</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>17</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,21,47.5,21</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,31,66,31</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<connection>
<GID>21</GID>
<name>N_in0</name></connection>
<intersection>61.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>61.5,16,61.5,31</points>
<intersection>16 5</intersection>
<intersection>31 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>47.5,16,61.5,16</points>
<intersection>47.5 6</intersection>
<intersection>61.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>47.5,16,47.5,23</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>16 5</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,22,66,22</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<connection>
<GID>23</GID>
<name>N_in0</name></connection>
<intersection>59 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>59,22,59,25.5</points>
<intersection>22 1</intersection>
<intersection>25.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>47.5,25.5,59,25.5</points>
<intersection>47.5 12</intersection>
<intersection>59 10</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>47.5,25.5,47.5,30</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>25.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,2,10.5,2</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-4,11,-4</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,2,36,2</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>34 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34,-6,34,2</points>
<intersection>-6 4</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>34,-6,44.5,-6</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>34 3</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,2,44.5,2</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-8,44.5,-8</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>40.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>40.5,-8,40.5,4</points>
<intersection>-8 1</intersection>
<intersection>4 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>40.5,4,44.5,4</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>40.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,3,58.5,3</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,2,72.5,2</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<connection>
<GID>41</GID>
<name>N_in0</name></connection>
<intersection>68 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>68,-2,68,2</points>
<intersection>-2 6</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>58.5,-2,68,-2</points>
<intersection>58.5 7</intersection>
<intersection>68 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>58.5,-5,58.5,-2</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-2 6</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-7,58.5,-7</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<connection>
<GID>42</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-3,69.5,-3</points>
<intersection>54.5 3</intersection>
<intersection>69.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54.5,-3,54.5,1</points>
<intersection>-3 1</intersection>
<intersection>1 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>54.5,1,58.5,1</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>54.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>69.5,-6,69.5,-3</points>
<intersection>-6 7</intersection>
<intersection>-6 7</intersection>
<intersection>-3 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>64.5,-6,72.5,-6</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<connection>
<GID>43</GID>
<name>N_in0</name></connection>
<intersection>69.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7.5,-83.5,-3,-83.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8,-149.5,-1,-149.5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8,-127,0.5,-127</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-8 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-8,-127,-8,-127</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>-127 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-149,81.5,-149</points>
<intersection>37.5 7</intersection>
<intersection>81.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>81.5,-149,81.5,-129</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>-149 1</intersection>
<intersection>-135.5 11</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>37.5,-149,37.5,-137.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>-149 1</intersection>
<intersection>-137.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>37.5,-137.5,43,-137.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>37.5 7</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>81.5,-135.5,82.5,-135.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>81.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,-137.5,54.5,-137.5</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>49.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49.5,-137.5,49.5,-129</points>
<intersection>-137.5 1</intersection>
<intersection>-129 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>49.5,-129,54,-129</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>49.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-127,54,-127</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<connection>
<GID>56</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-135.5,54,-132</points>
<intersection>-135.5 2</intersection>
<intersection>-132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-132,64.5,-132</points>
<intersection>54 0</intersection>
<intersection>64.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-135.5,54.5,-135.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>64.5,-132,64.5,-127</points>
<intersection>-132 1</intersection>
<intersection>-128 6</intersection>
<intersection>-127 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>64.5,-127,68,-127</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>64.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>60,-128,64.5,-128</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>64.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-137.5,64.5,-136.5</points>
<intersection>-137.5 2</intersection>
<intersection>-136.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-136.5,64.5,-136.5</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-137.5,68.5,-137.5</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-133.5,66,-129</points>
<intersection>-133.5 1</intersection>
<intersection>-129 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66,-133.5,75,-133.5</points>
<intersection>66 0</intersection>
<intersection>75 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66,-129,68,-129</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>66 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75,-137.5,75,-133.5</points>
<intersection>-137.5 4</intersection>
<intersection>-136.5 5</intersection>
<intersection>-133.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>75,-137.5,82.5,-137.5</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>75 3</intersection>
<intersection>75.5 6</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>74.5,-136.5,75,-136.5</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<intersection>75 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>75.5,-143,75.5,-137.5</points>
<connection>
<GID>62</GID>
<name>N_in3</name></connection>
<intersection>-137.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-131.5,74.5,-127</points>
<intersection>-131.5 2</intersection>
<intersection>-128 4</intersection>
<intersection>-127 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-127,81.5,-127</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection>
<intersection>75.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68.5,-131.5,74.5,-131.5</points>
<intersection>68.5 3</intersection>
<intersection>74.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>68.5,-135.5,68.5,-131.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>-131.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>74,-128,74.5,-128</points>
<connection>
<GID>57</GID>
<name>OUT</name></connection>
<intersection>74.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>75.5,-127,75.5,-122.5</points>
<connection>
<GID>61</GID>
<name>N_in2</name></connection>
<intersection>-127 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-81.5,77.5,-81.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>62.5 4</intersection>
<intersection>70 5</intersection>
<intersection>75.5 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>62.5,-82,62.5,-81.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>-81.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>70,-86.5,70,-81.5</points>
<connection>
<GID>22</GID>
<name>N_in3</name></connection>
<intersection>-81.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>75.5,-81.5,75.5,-78</points>
<intersection>-81.5 1</intersection>
<intersection>-78 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>56.5,-78,75.5,-78</points>
<intersection>56.5 8</intersection>
<intersection>75.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>56.5,-78,56.5,-75</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>-78 7</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-77,77.5,-77</points>
<intersection>54 5</intersection>
<intersection>67.5 8</intersection>
<intersection>70.5 4</intersection>
<intersection>77.5 7</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>70.5,-77,70.5,-68</points>
<connection>
<GID>18</GID>
<name>N_in2</name></connection>
<intersection>-77 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>54,-81,54,-77</points>
<intersection>-81 6</intersection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>54,-81,56.5,-81</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>54 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>77.5,-77,77.5,-74</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>-77 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>67.5,-77,67.5,-74</points>
<intersection>-77 1</intersection>
<intersection>-74 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>62.5,-74,67.5,-74</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>67.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-144,76.5,-144</points>
<connection>
<GID>62</GID>
<name>N_in1</name></connection>
<connection>
<GID>62</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-128,93,-126.5</points>
<intersection>-128 2</intersection>
<intersection>-126.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-126.5,99,-126.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-128,93,-128</points>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<intersection>93 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-138,93.5,-136.5</points>
<intersection>-138 1</intersection>
<intersection>-136.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-138,99,-138</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>88.5,-136.5,93.5,-136.5</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-137.5,110.5,-134</points>
<intersection>-137.5 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-137.5,115,-137.5</points>
<connection>
<GID>68</GID>
<name>N_in0</name></connection>
<intersection>105 5</intersection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96,-134,110.5,-134</points>
<intersection>96 4</intersection>
<intersection>110.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>96,-134,96,-128.5</points>
<intersection>-134 2</intersection>
<intersection>-128.5 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>105,-137.5,105,-137</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>-137.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>96,-128.5,99,-128.5</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<intersection>96 4</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-94,73.5,-94</points>
<intersection>34 4</intersection>
<intersection>73.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>73.5,-94,73.5,-72</points>
<intersection>-94 1</intersection>
<intersection>-83.5 7</intersection>
<intersection>-72 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>34,-94,34,-84</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>-94 1</intersection>
<intersection>-84 10</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>73.5,-72,77.5,-72</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>73.5 2</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>73.5,-83.5,77.5,-83.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>73.5 2</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>31.5,-84,34,-84</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>34 4</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-74,42.5,-74</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>31.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31.5,-78.5,31.5,-74</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>-74 1</intersection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-82,39,-78.5</points>
<intersection>-82 1</intersection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-82,44.5,-82</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-78.5,39,-78.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-84,44.5,-84</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>41 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>41,-84,41,-72</points>
<intersection>-84 1</intersection>
<intersection>-72 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>41,-72,42.5,-72</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>41 3</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-83,56.5,-83</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<connection>
<GID>15</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-73,56.5,-73</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-82.5,90.5,-82.5</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<connection>
<GID>26</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-73,86.5,-72</points>
<intersection>-73 2</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-72,90,-72</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,-73,86.5,-73</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-130.5,108.5,-126.5</points>
<intersection>-130.5 2</intersection>
<intersection>-126.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-126.5,114.5,-126.5</points>
<intersection>105 5</intersection>
<intersection>108.5 0</intersection>
<intersection>114.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-130.5,108.5,-130.5</points>
<intersection>99 6</intersection>
<intersection>108.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>114.5,-127.5,114.5,-126.5</points>
<connection>
<GID>67</GID>
<name>N_in0</name></connection>
<intersection>-126.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>105,-127.5,105,-126.5</points>
<connection>
<GID>65</GID>
<name>OUT</name></connection>
<intersection>-126.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>99,-136,99,-130.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>-130.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-76.5,108,-73</points>
<intersection>-76.5 4</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96,-73,109.5,-73</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<connection>
<GID>48</GID>
<name>N_in0</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>90.5,-76.5,108,-76.5</points>
<intersection>90.5 5</intersection>
<intersection>108 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>90.5,-80.5,90.5,-76.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-76.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96.5,-81.5,109,-81.5</points>
<connection>
<GID>52</GID>
<name>N_in0</name></connection>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>101 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>101,-81.5,101,-78</points>
<intersection>-81.5 1</intersection>
<intersection>-78 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>87.5,-78,101,-78</points>
<intersection>87.5 5</intersection>
<intersection>101 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>87.5,-78,87.5,-74</points>
<intersection>-78 4</intersection>
<intersection>-74 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>87.5,-74,90,-74</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>87.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-14.5,-195,-3.5,-195</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>-3.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-3.5,-195,-3.5,-195</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>-195 1</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-173.5,-2.5,-173.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-178.5,51.5,-178.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>31.5 3</intersection>
<intersection>35 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31.5,-181,31.5,-178.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>-178.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>35,-181,35,-178.5</points>
<intersection>-181 5</intersection>
<intersection>-178.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>35,-181,38,-181</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>35 4</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-180.5,66.5,-180.5</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<connection>
<GID>88</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-194.5,66.5,-194.5</points>
<connection>
<GID>86</GID>
<name>OUT</name></connection>
<connection>
<GID>89</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-14,-207.5,0,-207.5</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<connection>
<GID>82</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-192.5,46.5,-181</points>
<intersection>-192.5 1</intersection>
<intersection>-181 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-192.5,51.5,-192.5</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42,-181,46.5,-181</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-188.5,80.5,-181.5</points>
<intersection>-188.5 2</intersection>
<intersection>-184 1</intersection>
<intersection>-181.5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-184,95,-184</points>
<intersection>80.5 0</intersection>
<intersection>95 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66.5,-188.5,80.5,-188.5</points>
<intersection>66.5 3</intersection>
<intersection>80.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>66.5,-192.5,66.5,-188.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>-188.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>95,-184,95,-183</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>-184 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>72.5,-181.5,80.5,-181.5</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<intersection>77.5 8</intersection>
<intersection>80.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>77.5,-181.5,77.5,-172</points>
<connection>
<GID>92</GID>
<name>N_in2</name></connection>
<intersection>-181.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-193.5,79,-186.5</points>
<intersection>-193.5 1</intersection>
<intersection>-193.5 1</intersection>
<intersection>-186.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-193.5,95.5,-193.5</points>
<connection>
<GID>89</GID>
<name>OUT</name></connection>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>77.5 3</intersection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66.5,-186.5,79,-186.5</points>
<intersection>66.5 4</intersection>
<intersection>79 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77.5,-199.5,77.5,-193.5</points>
<connection>
<GID>94</GID>
<name>N_in3</name></connection>
<intersection>-193.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>66.5,-186.5,66.5,-182.5</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<intersection>-186.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-196,109.5,-194.5</points>
<intersection>-196 1</intersection>
<intersection>-194.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-196,118,-196</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101.5,-194.5,109.5,-194.5</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-182,108.5,-181</points>
<intersection>-182 2</intersection>
<intersection>-181 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-181,116.5,-181</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101,-182,108.5,-182</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-182,151,-181</points>
<connection>
<GID>104</GID>
<name>N_in3</name></connection>
<intersection>-182 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-182,151,-182</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<intersection>129.5 5</intersection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>129.5,-190,129.5,-182</points>
<intersection>-190 6</intersection>
<intersection>-182 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>113,-190,129.5,-190</points>
<intersection>113 7</intersection>
<intersection>129.5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>113,-194,113,-190</points>
<intersection>-194 8</intersection>
<intersection>-190 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>113,-194,118,-194</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>113 7</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-195,150.5,-195</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<connection>
<GID>106</GID>
<name>N_in0</name></connection>
<intersection>135.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>135.5,-195,135.5,-187.5</points>
<intersection>-195 1</intersection>
<intersection>-187.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>113,-187.5,135.5,-187.5</points>
<intersection>113 6</intersection>
<intersection>135.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>113,-187.5,113,-183</points>
<intersection>-187.5 5</intersection>
<intersection>-183 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>113,-183,116.5,-183</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>113 6</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-194.5,49,-180.5</points>
<intersection>-194.5 3</intersection>
<intersection>-187 4</intersection>
<intersection>-180.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-180.5,51.5,-180.5</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>49,-194.5,51.5,-194.5</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>44,-187,49,-187</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-211.5,63,-202</points>
<intersection>-211.5 1</intersection>
<intersection>-202 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-211.5,95.5,-211.5</points>
<intersection>63 0</intersection>
<intersection>88 4</intersection>
<intersection>95.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-202,63,-202</points>
<intersection>38.5 6</intersection>
<intersection>63 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>95.5,-211.5,95.5,-195.5</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>-211.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>88,-211.5,88,-181</points>
<intersection>-211.5 1</intersection>
<intersection>-181 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>88,-181,95,-181</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>88 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>38.5,-202,38.5,-187</points>
<intersection>-202 2</intersection>
<intersection>-187 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>31,-187,40,-187</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>38.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-196.5,42,-182.5</points>
<intersection>-196.5 3</intersection>
<intersection>-194.5 2</intersection>
<intersection>-182.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-182.5,51.5,-182.5</points>
<connection>
<GID>85</GID>
<name>IN_2</name></connection>
<intersection>42 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-194.5,42,-194.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>42 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>42,-196.5,51.5,-196.5</points>
<connection>
<GID>86</GID>
<name>IN_2</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-7.02185,0,303.987,-343.025</PageViewport></page 1>
<page 2>
<PageViewport>-7.02185,0,303.987,-343.025</PageViewport></page 2>
<page 3>
<PageViewport>-7.02185,0,303.987,-343.025</PageViewport></page 3>
<page 4>
<PageViewport>-7.02185,0,303.987,-343.025</PageViewport></page 4>
<page 5>
<PageViewport>-7.02185,0,303.987,-343.025</PageViewport></page 5>
<page 6>
<PageViewport>-7.02185,0,303.987,-343.025</PageViewport></page 6>
<page 7>
<PageViewport>-7.02185,0,303.987,-343.025</PageViewport></page 7>
<page 8>
<PageViewport>-7.02185,0,303.987,-343.025</PageViewport></page 8>
<page 9>
<PageViewport>-7.02185,0,303.987,-343.025</PageViewport></page 9></circuit>