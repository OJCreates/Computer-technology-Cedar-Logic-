<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>21.3029,30.2381,126.265,-83.8508</PageViewport>
<gate>
<ID>10</ID>
<type>DD_KEYPAD_HEX</type>
<position>19,-35</position>
<output>
<ID>OUT_0</ID>6 </output>
<output>
<ID>OUT_1</ID>5 </output>
<output>
<ID>OUT_2</ID>4 </output>
<output>
<ID>OUT_3</ID>3 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>12</ID>
<type>DE_TO</type>
<position>35,-32</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>13</ID>
<type>DE_TO</type>
<position>35,-34</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>14</ID>
<type>DE_TO</type>
<position>35,-36</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>15</ID>
<type>DE_TO</type>
<position>35,-38</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>17,-45.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>21</ID>
<type>DE_TO</type>
<position>26.5,-45.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_REGISTER4</type>
<position>66.5,-22</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>9 </input>
<input>
<ID>IN_3</ID>8 </input>
<input>
<ID>clear</ID>21 </input>
<input>
<ID>clock</ID>20 </input>
<input>
<ID>count_enable</ID>108 </input>
<input>
<ID>count_up</ID>109 </input>
<input>
<ID>load</ID>24 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_REGISTER4</type>
<position>90,-22</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>13 </input>
<input>
<ID>IN_3</ID>12 </input>
<input>
<ID>clear</ID>22 </input>
<input>
<ID>clock</ID>20 </input>
<input>
<ID>count_enable</ID>45 </input>
<input>
<ID>count_up</ID>41 </input>
<input>
<ID>load</ID>26 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_REGISTER4</type>
<position>114,-22</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>16 </input>
<input>
<ID>clear</ID>23 </input>
<input>
<ID>clock</ID>20 </input>
<input>
<ID>count_enable</ID>110 </input>
<input>
<ID>count_up</ID>111 </input>
<input>
<ID>load</ID>27 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>29</ID>
<type>DA_FROM</type>
<position>57.5,-20</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>51.5,-21</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>57.5,-22</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>51.5,-23</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>80.5,-20</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>75.5,-21</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>80.5,-22</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>75.5,-23</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>37</ID>
<type>DA_FROM</type>
<position>106,-20</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>38</ID>
<type>DA_FROM</type>
<position>101,-21</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>39</ID>
<type>DA_FROM</type>
<position>106,-22</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>40</ID>
<type>DA_FROM</type>
<position>101,-23</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>58.5,-31</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>44</ID>
<type>FF_GND</type>
<position>67.5,-28.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>46</ID>
<type>FF_GND</type>
<position>91,-28.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>FF_GND</type>
<position>115,-28.5</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>DA_FROM</type>
<position>56.5,-14</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L0</lparam></gate>
<gate>
<ID>54</ID>
<type>DA_FROM</type>
<position>81,-13.5</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L1</lparam></gate>
<gate>
<ID>55</ID>
<type>DA_FROM</type>
<position>104,-13.5</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L2</lparam></gate>
<gate>
<ID>77</ID>
<type>EE_VDD</type>
<position>90,-13</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>78</ID>
<type>EE_VDD</type>
<position>92,-11.5</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>108</ID>
<type>FF_GND</type>
<position>66.5,-8</position>
<output>
<ID>OUT_0</ID>108 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>109</ID>
<type>FF_GND</type>
<position>68.5,-7</position>
<output>
<ID>OUT_0</ID>109 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>110</ID>
<type>FF_GND</type>
<position>113.5,-11</position>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>111</ID>
<type>FF_GND</type>
<position>115.5,-10.5</position>
<output>
<ID>OUT_0</ID>111 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-32,33,-32</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-34,33,-34</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-36,33,-36</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-38,33,-38</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-45.5,24.5,-45.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<connection>
<GID>21</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-20,62.5,-20</points>
<connection>
<GID>23</GID>
<name>IN_3</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-21,62.5,-21</points>
<connection>
<GID>23</GID>
<name>IN_2</name></connection>
<connection>
<GID>30</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-22,62.5,-22</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<connection>
<GID>31</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-23,62.5,-23</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-20,86,-20</points>
<connection>
<GID>25</GID>
<name>IN_3</name></connection>
<connection>
<GID>33</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>77.5,-21,86,-21</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<connection>
<GID>34</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-22,86,-22</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<connection>
<GID>35</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>77.5,-23,86,-23</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-20,110,-20</points>
<connection>
<GID>27</GID>
<name>IN_3</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-21,110,-21</points>
<connection>
<GID>27</GID>
<name>IN_2</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-22,110,-22</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-23,110,-23</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-31,65.5,-26</points>
<connection>
<GID>23</GID>
<name>clock</name></connection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-31,113,-31</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection>
<intersection>89 3</intersection>
<intersection>113 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>89,-31,89,-26</points>
<connection>
<GID>25</GID>
<name>clock</name></connection>
<intersection>-31 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>113,-31,113,-26</points>
<connection>
<GID>27</GID>
<name>clock</name></connection>
<intersection>-31 1</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-27.5,67.5,-26</points>
<connection>
<GID>23</GID>
<name>clear</name></connection>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-27.5,91,-26</points>
<connection>
<GID>25</GID>
<name>clear</name></connection>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-27.5,115,-26</points>
<connection>
<GID>27</GID>
<name>clear</name></connection>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-17,65.5,-14</points>
<connection>
<GID>23</GID>
<name>load</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-14,65.5,-14</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-17,89,-13.5</points>
<connection>
<GID>25</GID>
<name>load</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-13.5,89,-13.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-17,113,-13.5</points>
<connection>
<GID>27</GID>
<name>load</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-13.5,113,-13.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-17,91,-14.5</points>
<connection>
<GID>25</GID>
<name>count_up</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>92,-14.5,92,-12.5</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>91,-14.5,92,-14.5</points>
<intersection>91 0</intersection>
<intersection>92 1</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-17,90,-14</points>
<connection>
<GID>25</GID>
<name>count_enable</name></connection>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-17,66.5,-9</points>
<connection>
<GID>23</GID>
<name>count_enable</name></connection>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-17,67.5,-12.5</points>
<connection>
<GID>23</GID>
<name>count_up</name></connection>
<intersection>-12.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>68.5,-12.5,68.5,-8</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>67.5,-12.5,68.5,-12.5</points>
<intersection>67.5 0</intersection>
<intersection>68.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-17,114,-14.5</points>
<connection>
<GID>27</GID>
<name>count_enable</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>113.5,-14.5,113.5,-12</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-14.5,114,-14.5</points>
<intersection>113.5 1</intersection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-17,115,-14</points>
<connection>
<GID>27</GID>
<name>count_up</name></connection>
<intersection>-14 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>115.5,-14,115.5,-11.5</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>115,-14,115.5,-14</points>
<intersection>115 0</intersection>
<intersection>115.5 1</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-93.7465,35,51.9961,-123.416</PageViewport>
<gate>
<ID>1</ID>
<type>DD_KEYPAD_HEX</type>
<position>12,-56.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<output>
<ID>OUT_1</ID>29 </output>
<output>
<ID>OUT_2</ID>28 </output>
<output>
<ID>OUT_3</ID>25 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>3</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>108,-57.5</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_2</ID>70 </input>
<input>
<ID>IN_3</ID>71 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>5</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>29,-57</position>
<input>
<ID>ENABLE_0</ID>79 </input>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>29 </input>
<input>
<ID>IN_2</ID>28 </input>
<input>
<ID>IN_3</ID>25 </input>
<output>
<ID>OUT_0</ID>72 </output>
<output>
<ID>OUT_1</ID>83 </output>
<output>
<ID>OUT_2</ID>70 </output>
<output>
<ID>OUT_3</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_REGISTER4</type>
<position>40.5,-36.5</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_2</ID>70 </input>
<input>
<ID>IN_3</ID>71 </input>
<output>
<ID>OUT_0</ID>40 </output>
<output>
<ID>OUT_1</ID>35 </output>
<output>
<ID>OUT_2</ID>39 </output>
<output>
<ID>OUT_3</ID>34 </output>
<input>
<ID>clear</ID>33 </input>
<input>
<ID>clock</ID>49 </input>
<input>
<ID>count_enable</ID>32 </input>
<input>
<ID>count_up</ID>31 </input>
<input>
<ID>load</ID>51 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>9</ID>
<type>FF_GND</type>
<position>41.5,-30.5</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>11</ID>
<type>FF_GND</type>
<position>40.5,-29</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>FF_GND</type>
<position>41.5,-41.5</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>47,-36</position>
<input>
<ID>ENABLE_0</ID>80 </input>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>35 </input>
<input>
<ID>IN_2</ID>39 </input>
<input>
<ID>IN_3</ID>34 </input>
<output>
<ID>OUT_0</ID>72 </output>
<output>
<ID>OUT_1</ID>83 </output>
<output>
<ID>OUT_2</ID>70 </output>
<output>
<ID>OUT_3</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>39.5,-42.5</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>20</ID>
<type>DE_TO</type>
<position>17,-69.5</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>10.5,-69.5</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>24</ID>
<type>BA_DECODER_2x4</type>
<position>24.5,-24</position>
<input>
<ID>ENABLE</ID>77 </input>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT_1</ID>51 </output>
<output>
<ID>OUT_2</ID>73 </output>
<output>
<ID>OUT_3</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>DD_KEYPAD_HEX</type>
<position>13.5,-23.5</position>
<output>
<ID>OUT_0</ID>52 </output>
<output>
<ID>OUT_1</ID>53 </output>
<output>
<ID>OUT_2</ID>75 </output>
<output>
<ID>OUT_3</ID>76 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_REGISTER4</type>
<position>62.5,-36.5</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_2</ID>70 </input>
<input>
<ID>IN_3</ID>71 </input>
<output>
<ID>OUT_0</ID>60 </output>
<output>
<ID>OUT_1</ID>58 </output>
<output>
<ID>OUT_2</ID>59 </output>
<output>
<ID>OUT_3</ID>57 </output>
<input>
<ID>clear</ID>56 </input>
<input>
<ID>clock</ID>61 </input>
<input>
<ID>count_enable</ID>55 </input>
<input>
<ID>count_up</ID>54 </input>
<input>
<ID>load</ID>73 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>41</ID>
<type>FF_GND</type>
<position>63.5,-30.5</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>43</ID>
<type>FF_GND</type>
<position>62.5,-29</position>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>45</ID>
<type>FF_GND</type>
<position>63.5,-41.5</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>47</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>69,-36</position>
<input>
<ID>ENABLE_0</ID>81 </input>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>57 </input>
<output>
<ID>OUT_0</ID>72 </output>
<output>
<ID>OUT_1</ID>83 </output>
<output>
<ID>OUT_2</ID>70 </output>
<output>
<ID>OUT_3</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>48</ID>
<type>DA_FROM</type>
<position>61.5,-42.5</position>
<input>
<ID>IN_0</ID>61 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_REGISTER4</type>
<position>90,-36.5</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_2</ID>70 </input>
<input>
<ID>IN_3</ID>71 </input>
<output>
<ID>OUT_0</ID>68 </output>
<output>
<ID>OUT_1</ID>66 </output>
<output>
<ID>OUT_2</ID>67 </output>
<output>
<ID>OUT_3</ID>65 </output>
<input>
<ID>clear</ID>64 </input>
<input>
<ID>clock</ID>69 </input>
<input>
<ID>count_enable</ID>63 </input>
<input>
<ID>count_up</ID>62 </input>
<input>
<ID>load</ID>74 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>52</ID>
<type>FF_GND</type>
<position>91,-30.5</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>53</ID>
<type>FF_GND</type>
<position>90,-29</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>FF_GND</type>
<position>91,-41.5</position>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>57</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>96.5,-36</position>
<input>
<ID>ENABLE_0</ID>82 </input>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>66 </input>
<input>
<ID>IN_2</ID>67 </input>
<input>
<ID>IN_3</ID>65 </input>
<output>
<ID>OUT_0</ID>72 </output>
<output>
<ID>OUT_1</ID>83 </output>
<output>
<ID>OUT_2</ID>70 </output>
<output>
<ID>OUT_3</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>89,-42.5</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>59</ID>
<type>BA_DECODER_2x4</type>
<position>25.5,-17.5</position>
<input>
<ID>ENABLE</ID>78 </input>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT_0</ID>79 </output>
<output>
<ID>OUT_1</ID>80 </output>
<output>
<ID>OUT_2</ID>81 </output>
<output>
<ID>OUT_3</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>EE_VDD</type>
<position>20,-16</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>61</ID>
<type>EE_VDD</type>
<position>19.5,-23.5</position>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-53.5,27,-53.5</points>
<connection>
<GID>1</GID>
<name>OUT_3</name></connection>
<intersection>27 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27,-55.5,27,-53.5</points>
<connection>
<GID>5</GID>
<name>IN_3</name></connection>
<intersection>-53.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-56.5,22,-55.5</points>
<intersection>-56.5 1</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-56.5,27,-56.5</points>
<connection>
<GID>5</GID>
<name>IN_2</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-55.5,22,-55.5</points>
<connection>
<GID>1</GID>
<name>OUT_2</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-57.5,27,-57.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<connection>
<GID>1</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-59.5,22,-58.5</points>
<intersection>-59.5 2</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-58.5,27,-58.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-59.5,22,-59.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>41.5,-31.5,41.5,-31.5</points>
<connection>
<GID>7</GID>
<name>count_up</name></connection>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-31.5,40.5,-30</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<connection>
<GID>7</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>41.5,-40.5,41.5,-40.5</points>
<connection>
<GID>7</GID>
<name>clear</name></connection>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>44.5,-34.5,45,-34.5</points>
<connection>
<GID>17</GID>
<name>IN_3</name></connection>
<connection>
<GID>7</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>44.5,-36.5,45,-36.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<connection>
<GID>7</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>44.5,-35.5,45,-35.5</points>
<connection>
<GID>17</GID>
<name>IN_2</name></connection>
<connection>
<GID>7</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>44.5,-37.5,45,-37.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>39.5,-40.5,39.5,-40.5</points>
<connection>
<GID>7</GID>
<name>clock</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,-69.5,15,-69.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-31.5,39.5,-24.5</points>
<connection>
<GID>7</GID>
<name>load</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-24.5,39.5,-24.5</points>
<connection>
<GID>24</GID>
<name>OUT_1</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-26.5,20,-25.5</points>
<intersection>-26.5 2</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-25.5,21.5,-25.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-26.5,20,-26.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,-24.5,21.5,-24.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<connection>
<GID>26</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>63.5,-31.5,63.5,-31.5</points>
<connection>
<GID>28</GID>
<name>count_up</name></connection>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-31.5,62.5,-30</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<connection>
<GID>28</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>63.5,-40.5,63.5,-40.5</points>
<connection>
<GID>28</GID>
<name>clear</name></connection>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>66.5,-34.5,67,-34.5</points>
<connection>
<GID>47</GID>
<name>IN_3</name></connection>
<connection>
<GID>28</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>66.5,-36.5,67,-36.5</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<connection>
<GID>28</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>66.5,-35.5,67,-35.5</points>
<connection>
<GID>47</GID>
<name>IN_2</name></connection>
<connection>
<GID>28</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>66.5,-37.5,67,-37.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>61.5,-40.5,61.5,-40.5</points>
<connection>
<GID>28</GID>
<name>clock</name></connection>
<connection>
<GID>48</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>91,-31.5,91,-31.5</points>
<connection>
<GID>50</GID>
<name>count_up</name></connection>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-31.5,90,-30</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<connection>
<GID>50</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>91,-40.5,91,-40.5</points>
<connection>
<GID>50</GID>
<name>clear</name></connection>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-34.5,94.5,-34.5</points>
<connection>
<GID>57</GID>
<name>IN_3</name></connection>
<connection>
<GID>50</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-36.5,94.5,-36.5</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<connection>
<GID>50</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-35.5,94.5,-35.5</points>
<connection>
<GID>57</GID>
<name>IN_2</name></connection>
<connection>
<GID>50</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-37.5,94.5,-37.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>89,-40.5,89,-40.5</points>
<connection>
<GID>50</GID>
<name>clock</name></connection>
<connection>
<GID>58</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-56.5,105,-56.5</points>
<connection>
<GID>5</GID>
<name>OUT_2</name></connection>
<connection>
<GID>3</GID>
<name>IN_2</name></connection>
<intersection>34.5 8</intersection>
<intersection>51 12</intersection>
<intersection>56.5 13</intersection>
<intersection>74 20</intersection>
<intersection>84 21</intersection>
<intersection>100.5 19</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>34.5,-56.5,34.5,-35.5</points>
<intersection>-56.5 1</intersection>
<intersection>-35.5 25</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>51,-56.5,51,-35.5</points>
<intersection>-56.5 1</intersection>
<intersection>-35.5 16</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>56.5,-56.5,56.5,-35.5</points>
<intersection>-56.5 1</intersection>
<intersection>-35.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>56.5,-35.5,58.5,-35.5</points>
<connection>
<GID>28</GID>
<name>IN_2</name></connection>
<intersection>56.5 13</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>49,-35.5,51,-35.5</points>
<connection>
<GID>17</GID>
<name>OUT_2</name></connection>
<intersection>51 12</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>100.5,-56.5,100.5,-35.5</points>
<intersection>-56.5 1</intersection>
<intersection>-35.5 24</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>74,-56.5,74,-35.5</points>
<intersection>-56.5 1</intersection>
<intersection>-35.5 22</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>84,-56.5,84,-35.5</points>
<intersection>-56.5 1</intersection>
<intersection>-35.5 23</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>71,-35.5,74,-35.5</points>
<connection>
<GID>47</GID>
<name>OUT_2</name></connection>
<intersection>74 20</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>84,-35.5,86,-35.5</points>
<connection>
<GID>50</GID>
<name>IN_2</name></connection>
<intersection>84 21</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>98.5,-35.5,100.5,-35.5</points>
<connection>
<GID>57</GID>
<name>OUT_2</name></connection>
<intersection>100.5 19</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>34.5,-35.5,36.5,-35.5</points>
<connection>
<GID>7</GID>
<name>IN_2</name></connection>
<intersection>34.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-55.5,105,-55.5</points>
<connection>
<GID>5</GID>
<name>OUT_3</name></connection>
<connection>
<GID>3</GID>
<name>IN_3</name></connection>
<intersection>33 9</intersection>
<intersection>51.5 13</intersection>
<intersection>55 14</intersection>
<intersection>75 23</intersection>
<intersection>83 24</intersection>
<intersection>102 22</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>33,-55.5,33,-34.5</points>
<intersection>-55.5 1</intersection>
<intersection>-34.5 29</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>51.5,-55.5,51.5,-34.5</points>
<intersection>-55.5 1</intersection>
<intersection>-34.5 28</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>55,-55.5,55,-34.5</points>
<intersection>-55.5 1</intersection>
<intersection>-34.5 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>55,-34.5,58.5,-34.5</points>
<connection>
<GID>28</GID>
<name>IN_3</name></connection>
<intersection>55 14</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>102,-55.5,102,-34.5</points>
<intersection>-55.5 1</intersection>
<intersection>-34.5 27</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>75,-55.5,75,-34.5</points>
<intersection>-55.5 1</intersection>
<intersection>-34.5 25</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>83,-55.5,83,-34.5</points>
<intersection>-55.5 1</intersection>
<intersection>-34.5 26</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>71,-34.5,75,-34.5</points>
<connection>
<GID>47</GID>
<name>OUT_3</name></connection>
<intersection>75 23</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>83,-34.5,86,-34.5</points>
<connection>
<GID>50</GID>
<name>IN_3</name></connection>
<intersection>83 24</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>98.5,-34.5,102,-34.5</points>
<connection>
<GID>57</GID>
<name>OUT_3</name></connection>
<intersection>102 22</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>49,-34.5,51.5,-34.5</points>
<connection>
<GID>17</GID>
<name>OUT_3</name></connection>
<intersection>51.5 13</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>33,-34.5,36.5,-34.5</points>
<connection>
<GID>7</GID>
<name>IN_3</name></connection>
<intersection>33 9</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-58.5,105,-58.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>36.5 4</intersection>
<intersection>49 6</intersection>
<intersection>58.5 10</intersection>
<intersection>71 9</intersection>
<intersection>86 14</intersection>
<intersection>98.5 13</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>36.5,-58.5,36.5,-37.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>49,-58.5,49,-37.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>71,-58.5,71,-37.5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>58.5,-58.5,58.5,-37.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>98.5,-58.5,98.5,-37.5</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>86,-58.5,86,-37.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>-58.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-31.5,61.5,-23.5</points>
<connection>
<GID>28</GID>
<name>load</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-23.5,61.5,-23.5</points>
<connection>
<GID>24</GID>
<name>OUT_2</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-31.5,89,-22.5</points>
<connection>
<GID>50</GID>
<name>load</name></connection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-22.5,89,-22.5</points>
<connection>
<GID>24</GID>
<name>OUT_3</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-22.5,21,-19</points>
<intersection>-22.5 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-22.5,21,-22.5</points>
<connection>
<GID>26</GID>
<name>OUT_2</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-19,22.5,-19</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-20.5,20,-18</points>
<intersection>-20.5 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-20.5,20,-20.5</points>
<connection>
<GID>26</GID>
<name>OUT_3</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,-18,22.5,-18</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-23.5,21.5,-22.5</points>
<connection>
<GID>24</GID>
<name>ENABLE</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-23.5,21.5,-23.5</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,-16,22.5,-16</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<connection>
<GID>59</GID>
<name>ENABLE</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-54,29,-19</points>
<connection>
<GID>5</GID>
<name>ENABLE_0</name></connection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-19,29,-19</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-33,47,-18</points>
<connection>
<GID>17</GID>
<name>ENABLE_0</name></connection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-18,47,-18</points>
<connection>
<GID>59</GID>
<name>OUT_1</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-33,69,-17</points>
<connection>
<GID>47</GID>
<name>ENABLE_0</name></connection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-17,69,-17</points>
<connection>
<GID>59</GID>
<name>OUT_2</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-33,96.5,-16</points>
<connection>
<GID>57</GID>
<name>ENABLE_0</name></connection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-16,96.5,-16</points>
<connection>
<GID>59</GID>
<name>OUT_3</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-57.5,105,-57.5</points>
<connection>
<GID>5</GID>
<name>OUT_1</name></connection>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>35.5 7</intersection>
<intersection>50 12</intersection>
<intersection>57.5 13</intersection>
<intersection>72.5 20</intersection>
<intersection>85 21</intersection>
<intersection>99.5 19</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>35.5,-57.5,35.5,-36.5</points>
<intersection>-57.5 1</intersection>
<intersection>-36.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>35.5,-36.5,36.5,-36.5</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>35.5 7</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>50,-57.5,50,-36.5</points>
<intersection>-57.5 1</intersection>
<intersection>-36.5 16</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>57.5,-57.5,57.5,-36.5</points>
<intersection>-57.5 1</intersection>
<intersection>-36.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>57.5,-36.5,58.5,-36.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>57.5 13</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>49,-36.5,50,-36.5</points>
<connection>
<GID>17</GID>
<name>OUT_1</name></connection>
<intersection>50 12</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>99.5,-57.5,99.5,-36.5</points>
<intersection>-57.5 1</intersection>
<intersection>-36.5 24</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>72.5,-57.5,72.5,-36.5</points>
<intersection>-57.5 1</intersection>
<intersection>-36.5 22</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>85,-57.5,85,-36.5</points>
<intersection>-57.5 1</intersection>
<intersection>-36.5 23</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>71,-36.5,72.5,-36.5</points>
<connection>
<GID>47</GID>
<name>OUT_1</name></connection>
<intersection>72.5 20</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>85,-36.5,86,-36.5</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>85 21</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>98.5,-36.5,99.5,-36.5</points>
<connection>
<GID>57</GID>
<name>OUT_1</name></connection>
<intersection>99.5 19</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>14.0898,40.5941,159.832,-117.822</PageViewport>
<gate>
<ID>62</ID>
<type>DD_KEYPAD_HEX</type>
<position>19,-21.5</position>
<output>
<ID>OUT_0</ID>91 </output>
<output>
<ID>OUT_1</ID>89 </output>
<output>
<ID>OUT_2</ID>86 </output>
<output>
<ID>OUT_3</ID>84 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 4</lparam></gate>
<gate>
<ID>64</ID>
<type>BA_DECODER_2x4</type>
<position>33,-14</position>
<input>
<ID>ENABLE</ID>85 </input>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT_0</ID>132 </output>
<output>
<ID>OUT_1</ID>131 </output>
<output>
<ID>OUT_2</ID>172 </output>
<output>
<ID>OUT_3</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>EE_VDD</type>
<position>27.5,-12.5</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>67</ID>
<type>BA_DECODER_2x4</type>
<position>30.5,-22</position>
<input>
<ID>ENABLE</ID>87 </input>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT_1</ID>112 </output>
<output>
<ID>OUT_2</ID>171 </output>
<output>
<ID>OUT_3</ID>173 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>EE_VDD</type>
<position>24.5,-21.5</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>75</ID>
<type>DD_KEYPAD_HEX</type>
<position>19.5,-55</position>
<output>
<ID>OUT_0</ID>95 </output>
<output>
<ID>OUT_1</ID>94 </output>
<output>
<ID>OUT_2</ID>93 </output>
<output>
<ID>OUT_3</ID>92 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>81</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>32,-55.5</position>
<input>
<ID>ENABLE_0</ID>132 </input>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>94 </input>
<input>
<ID>IN_2</ID>93 </input>
<input>
<ID>IN_3</ID>92 </input>
<output>
<ID>OUT_0</ID>103 </output>
<output>
<ID>OUT_1</ID>102 </output>
<output>
<ID>OUT_2</ID>101 </output>
<output>
<ID>OUT_3</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>85</ID>
<type>DE_TO</type>
<position>27,-71.5</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_TOGGLE</type>
<position>16.5,-71.5</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>96</ID>
<type>DE_TO</type>
<position>36.5,-54</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>97</ID>
<type>DE_TO</type>
<position>47,-55</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>98</ID>
<type>DE_TO</type>
<position>58.5,-56</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>99</ID>
<type>DE_TO</type>
<position>68.5,-57.5</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>101</ID>
<type>DA_FROM</type>
<position>50.5,-48.5</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>103</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>88,-50.5</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>106 </input>
<input>
<ID>IN_2</ID>105 </input>
<input>
<ID>IN_3</ID>104 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>104</ID>
<type>DA_FROM</type>
<position>59.5,-49.5</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>105</ID>
<type>DA_FROM</type>
<position>68.5,-50.5</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>106</ID>
<type>DA_FROM</type>
<position>77,-51.5</position>
<input>
<ID>IN_0</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_REGISTER4</type>
<position>47.5,-30</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>119 </input>
<input>
<ID>IN_2</ID>121 </input>
<input>
<ID>IN_3</ID>122 </input>
<output>
<ID>OUT_0</ID>126 </output>
<output>
<ID>OUT_1</ID>125 </output>
<output>
<ID>OUT_2</ID>124 </output>
<output>
<ID>OUT_3</ID>123 </output>
<input>
<ID>clear</ID>116 </input>
<input>
<ID>clock</ID>115 </input>
<input>
<ID>count_enable</ID>189 </input>
<input>
<ID>count_up</ID>188 </input>
<input>
<ID>load</ID>112 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>118</ID>
<type>DA_FROM</type>
<position>46.5,-36.5</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>119</ID>
<type>FF_GND</type>
<position>48.5,-35</position>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>120</ID>
<type>DA_FROM</type>
<position>41,-34.5</position>
<input>
<ID>IN_0</ID>118 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>121</ID>
<type>DA_FROM</type>
<position>37.5,-34.5</position>
<input>
<ID>IN_0</ID>119 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>122</ID>
<type>DA_FROM</type>
<position>34.5,-34.5</position>
<input>
<ID>IN_0</ID>121 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>123</ID>
<type>DA_FROM</type>
<position>31,-34.5</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>124</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>56,-29.5</position>
<input>
<ID>ENABLE_0</ID>131 </input>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>125 </input>
<input>
<ID>IN_2</ID>124 </input>
<input>
<ID>IN_3</ID>123 </input>
<output>
<ID>OUT_0</ID>130 </output>
<output>
<ID>OUT_1</ID>129 </output>
<output>
<ID>OUT_2</ID>128 </output>
<output>
<ID>OUT_3</ID>127 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>125</ID>
<type>DE_TO</type>
<position>69.5,-32.5</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>126</ID>
<type>DE_TO</type>
<position>66,-32.5</position>
<input>
<ID>IN_0</ID>128 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>127</ID>
<type>DE_TO</type>
<position>63,-32.5</position>
<input>
<ID>IN_0</ID>129 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>128</ID>
<type>DE_TO</type>
<position>60.5,-33</position>
<input>
<ID>IN_0</ID>130 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_REGISTER4</type>
<position>158,-22</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>140 </input>
<input>
<ID>IN_2</ID>150 </input>
<input>
<ID>IN_3</ID>149 </input>
<output>
<ID>OUT_0</ID>144 </output>
<output>
<ID>OUT_1</ID>143 </output>
<output>
<ID>OUT_2</ID>142 </output>
<output>
<ID>OUT_3</ID>141 </output>
<input>
<ID>clear</ID>138 </input>
<input>
<ID>clock</ID>137 </input>
<input>
<ID>count_enable</ID>182 </input>
<input>
<ID>count_up</ID>181 </input>
<input>
<ID>load</ID>173 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>141</ID>
<type>DA_FROM</type>
<position>157,-28.5</position>
<input>
<ID>IN_0</ID>137 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>142</ID>
<type>FF_GND</type>
<position>159,-27</position>
<output>
<ID>OUT_0</ID>138 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>143</ID>
<type>DA_FROM</type>
<position>151.5,-26.5</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>144</ID>
<type>DA_FROM</type>
<position>148,-26.5</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>145</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>166.5,-21.5</position>
<input>
<ID>ENABLE_0</ID>153 </input>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>143 </input>
<input>
<ID>IN_2</ID>142 </input>
<input>
<ID>IN_3</ID>141 </input>
<output>
<ID>OUT_0</ID>148 </output>
<output>
<ID>OUT_1</ID>147 </output>
<output>
<ID>OUT_2</ID>146 </output>
<output>
<ID>OUT_3</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>146</ID>
<type>DE_TO</type>
<position>180,-24.5</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>147</ID>
<type>DE_TO</type>
<position>176.5,-24.5</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>148</ID>
<type>DE_TO</type>
<position>173.5,-24.5</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>149</ID>
<type>DE_TO</type>
<position>171,-25</position>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>150</ID>
<type>DA_FROM</type>
<position>144.5,-26.5</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>151</ID>
<type>DA_FROM</type>
<position>140.5,-26.5</position>
<input>
<ID>IN_0</ID>149 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_REGISTER4</type>
<position>95.5,-27</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>158 </input>
<input>
<ID>IN_2</ID>168 </input>
<input>
<ID>IN_3</ID>167 </input>
<output>
<ID>OUT_0</ID>162 </output>
<output>
<ID>OUT_1</ID>161 </output>
<output>
<ID>OUT_2</ID>160 </output>
<output>
<ID>OUT_3</ID>159 </output>
<input>
<ID>clear</ID>156 </input>
<input>
<ID>clock</ID>155 </input>
<input>
<ID>count_enable</ID>187 </input>
<input>
<ID>count_up</ID>186 </input>
<input>
<ID>load</ID>171 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>156</ID>
<type>DA_FROM</type>
<position>94.5,-33.5</position>
<input>
<ID>IN_0</ID>155 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>157</ID>
<type>FF_GND</type>
<position>96.5,-32</position>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>158</ID>
<type>DA_FROM</type>
<position>89,-31.5</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>159</ID>
<type>DA_FROM</type>
<position>85.5,-31.5</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>160</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>104,-26.5</position>
<input>
<ID>ENABLE_0</ID>172 </input>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>161 </input>
<input>
<ID>IN_2</ID>160 </input>
<input>
<ID>IN_3</ID>159 </input>
<output>
<ID>OUT_0</ID>166 </output>
<output>
<ID>OUT_1</ID>165 </output>
<output>
<ID>OUT_2</ID>164 </output>
<output>
<ID>OUT_3</ID>163 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>161</ID>
<type>DE_TO</type>
<position>117.5,-29.5</position>
<input>
<ID>IN_0</ID>163 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>162</ID>
<type>DE_TO</type>
<position>114,-29.5</position>
<input>
<ID>IN_0</ID>164 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>163</ID>
<type>DE_TO</type>
<position>111,-29.5</position>
<input>
<ID>IN_0</ID>165 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 1</lparam></gate>
<gate>
<ID>164</ID>
<type>DE_TO</type>
<position>108.5,-30</position>
<input>
<ID>IN_0</ID>166 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Bus 0</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_FROM</type>
<position>82,-31.5</position>
<input>
<ID>IN_0</ID>168 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 2</lparam></gate>
<gate>
<ID>166</ID>
<type>DA_FROM</type>
<position>78,-31.5</position>
<input>
<ID>IN_0</ID>167 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Bus 3</lparam></gate>
<gate>
<ID>178</ID>
<type>FF_GND</type>
<position>159,-15</position>
<output>
<ID>OUT_0</ID>181 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>179</ID>
<type>FF_GND</type>
<position>158,-14.5</position>
<output>
<ID>OUT_0</ID>182 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>183</ID>
<type>FF_GND</type>
<position>95.5,-20.5</position>
<output>
<ID>OUT_0</ID>187 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>184</ID>
<type>FF_GND</type>
<position>96.5,-18.5</position>
<output>
<ID>OUT_0</ID>186 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>185</ID>
<type>FF_GND</type>
<position>47.5,-23.5</position>
<output>
<ID>OUT_0</ID>189 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>186</ID>
<type>FF_GND</type>
<position>48.5,-20.5</position>
<output>
<ID>OUT_0</ID>188 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-18.5,27,-14.5</points>
<intersection>-18.5 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-14.5,30,-14.5</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-18.5,27,-18.5</points>
<connection>
<GID>62</GID>
<name>OUT_3</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-12.5,30,-12.5</points>
<connection>
<GID>64</GID>
<name>ENABLE</name></connection>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-19.5,27.5,-15.5</points>
<intersection>-19.5 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-15.5,30,-15.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-19.5,27.5,-19.5</points>
<intersection>24 3</intersection>
<intersection>27.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24,-20.5,24,-19.5</points>
<connection>
<GID>62</GID>
<name>OUT_2</name></connection>
<intersection>-19.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-21.5,26.5,-20.5</points>
<intersection>-21.5 2</intersection>
<intersection>-20.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-21.5,26.5,-21.5</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26.5,-20.5,27.5,-20.5</points>
<connection>
<GID>67</GID>
<name>ENABLE</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-22.5,27.5,-22.5</points>
<connection>
<GID>62</GID>
<name>OUT_1</name></connection>
<connection>
<GID>67</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-24.5,25.5,-23.5</points>
<intersection>-24.5 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-23.5,27.5,-23.5</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-24.5,25.5,-24.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-54,30,-52</points>
<connection>
<GID>81</GID>
<name>IN_3</name></connection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-52,30,-52</points>
<connection>
<GID>75</GID>
<name>OUT_3</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-55,27,-54</points>
<intersection>-55 1</intersection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-55,30,-55</points>
<connection>
<GID>81</GID>
<name>IN_2</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-54,27,-54</points>
<connection>
<GID>75</GID>
<name>OUT_2</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-56,30,-56</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<connection>
<GID>75</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-58,27,-57</points>
<intersection>-58 2</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-57,30,-57</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-58,27,-58</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,-71.5,25,-71.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-54,34.5,-54</points>
<connection>
<GID>81</GID>
<name>OUT_3</name></connection>
<connection>
<GID>96</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-55,45,-55</points>
<connection>
<GID>81</GID>
<name>OUT_2</name></connection>
<connection>
<GID>97</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-56,56.5,-56</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<connection>
<GID>81</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-57.5,50,-57</points>
<intersection>-57.5 2</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-57,50,-57</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-57.5,66.5,-57.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,-48.5,85,-48.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<connection>
<GID>103</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61.5,-49.5,85,-49.5</points>
<connection>
<GID>103</GID>
<name>IN_2</name></connection>
<connection>
<GID>104</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-50.5,85,-50.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>85 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>85,-50.5,85,-50.5</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>-50.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79,-51.5,85,-51.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>85 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>85,-51.5,85,-51.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-25,46.5,-22.5</points>
<connection>
<GID>113</GID>
<name>load</name></connection>
<intersection>-22.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>33.5,-22.5,46.5,-22.5</points>
<connection>
<GID>67</GID>
<name>OUT_1</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-34.5,46.5,-34</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<connection>
<GID>113</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>48.5,-34,48.5,-34</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<connection>
<GID>113</GID>
<name>clear</name></connection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-32.5,41,-31</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-31,43.5,-31</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-32.5,37.5,-30</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-30,43.5,-30</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-32.5,34.5,-29</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-29,43.5,-29</points>
<connection>
<GID>113</GID>
<name>IN_2</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-32.5,31,-28</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-28,43.5,-28</points>
<connection>
<GID>113</GID>
<name>IN_3</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-28,54,-28</points>
<connection>
<GID>124</GID>
<name>IN_3</name></connection>
<connection>
<GID>113</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-29,54,-29</points>
<connection>
<GID>124</GID>
<name>IN_2</name></connection>
<connection>
<GID>113</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-30,54,-30</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<connection>
<GID>113</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-31,54,-31</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-30.5,69.5,-28</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-28,69.5,-28</points>
<connection>
<GID>124</GID>
<name>OUT_3</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-30.5,66,-29</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-29,66,-29</points>
<connection>
<GID>124</GID>
<name>OUT_2</name></connection>
<intersection>66 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-30.5,63,-30</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-30,63,-30</points>
<connection>
<GID>124</GID>
<name>OUT_1</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58,-31,60.5,-31</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-26.5,56,-14.5</points>
<connection>
<GID>124</GID>
<name>ENABLE_0</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-14.5,56,-14.5</points>
<connection>
<GID>64</GID>
<name>OUT_1</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-52.5,39.5,-15.5</points>
<intersection>-52.5 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-15.5,39.5,-15.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-52.5,39.5,-52.5</points>
<connection>
<GID>81</GID>
<name>ENABLE_0</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-26.5,157,-26</points>
<connection>
<GID>140</GID>
<name>clock</name></connection>
<connection>
<GID>141</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-26,159,-26</points>
<connection>
<GID>140</GID>
<name>clear</name></connection>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,-24.5,151.5,-23</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151.5,-23,154,-23</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>151.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-24.5,148,-22</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148,-22,154,-22</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-20,164.5,-20</points>
<connection>
<GID>140</GID>
<name>OUT_3</name></connection>
<connection>
<GID>145</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-21,164.5,-21</points>
<connection>
<GID>140</GID>
<name>OUT_2</name></connection>
<connection>
<GID>145</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-22,164.5,-22</points>
<connection>
<GID>140</GID>
<name>OUT_1</name></connection>
<connection>
<GID>145</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-23,164.5,-23</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<connection>
<GID>145</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180,-22.5,180,-20</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,-20,180,-20</points>
<connection>
<GID>145</GID>
<name>OUT_3</name></connection>
<intersection>180 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176.5,-22.5,176.5,-21</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,-21,176.5,-21</points>
<connection>
<GID>145</GID>
<name>OUT_2</name></connection>
<intersection>176.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173.5,-22.5,173.5,-22</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,-22,173.5,-22</points>
<connection>
<GID>145</GID>
<name>OUT_1</name></connection>
<intersection>173.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>168.5,-23,171,-23</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<connection>
<GID>145</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>140.5,-20,154,-20</points>
<connection>
<GID>140</GID>
<name>IN_3</name></connection>
<intersection>140.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>140.5,-24.5,140.5,-20</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-24.5,144.5,-21</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144.5,-21,154,-21</points>
<connection>
<GID>140</GID>
<name>IN_2</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,-18.5,166.5,-12.5</points>
<connection>
<GID>145</GID>
<name>ENABLE_0</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-12.5,166.5,-12.5</points>
<connection>
<GID>64</GID>
<name>OUT_3</name></connection>
<intersection>166.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,-31.5,94.5,-31</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<connection>
<GID>155</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-31,96.5,-31</points>
<connection>
<GID>155</GID>
<name>clear</name></connection>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-29.5,89,-28</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89,-28,91.5,-28</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-29.5,85.5,-27</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-27,91.5,-27</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99.5,-25,102,-25</points>
<connection>
<GID>155</GID>
<name>OUT_3</name></connection>
<connection>
<GID>160</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99.5,-26,102,-26</points>
<connection>
<GID>155</GID>
<name>OUT_2</name></connection>
<connection>
<GID>160</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99.5,-27,102,-27</points>
<connection>
<GID>155</GID>
<name>OUT_1</name></connection>
<connection>
<GID>160</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99.5,-28,102,-28</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<connection>
<GID>160</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-27.5,117.5,-25</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-25,117.5,-25</points>
<connection>
<GID>160</GID>
<name>OUT_3</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-27.5,114,-26</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-26,114,-26</points>
<connection>
<GID>160</GID>
<name>OUT_2</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-27.5,111,-27</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-27,111,-27</points>
<connection>
<GID>160</GID>
<name>OUT_1</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106,-28,108.5,-28</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-25,91.5,-25</points>
<connection>
<GID>155</GID>
<name>IN_3</name></connection>
<intersection>78 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78,-29.5,78,-25</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>-25 1</intersection></vsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-29.5,82,-26</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-26,91.5,-26</points>
<connection>
<GID>155</GID>
<name>IN_2</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,-22,94.5,-21.5</points>
<connection>
<GID>155</GID>
<name>load</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-21.5,94.5,-21.5</points>
<connection>
<GID>67</GID>
<name>OUT_2</name></connection>
<intersection>94.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-23.5,104,-13.5</points>
<connection>
<GID>160</GID>
<name>ENABLE_0</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-13.5,104,-13.5</points>
<connection>
<GID>64</GID>
<name>OUT_2</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-17,157,-15.5</points>
<connection>
<GID>140</GID>
<name>load</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-15.5,157,-15.5</points>
<intersection>33.5 2</intersection>
<intersection>157 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>33.5,-20.5,33.5,-15.5</points>
<connection>
<GID>67</GID>
<name>OUT_3</name></connection>
<intersection>-15.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-17,159,-16</points>
<connection>
<GID>140</GID>
<name>count_up</name></connection>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,-17,158,-15.5</points>
<connection>
<GID>140</GID>
<name>count_enable</name></connection>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-22,96.5,-19.5</points>
<connection>
<GID>155</GID>
<name>count_up</name></connection>
<connection>
<GID>184</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-22,95.5,-21.5</points>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection>
<connection>
<GID>155</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-25,48.5,-21.5</points>
<connection>
<GID>113</GID>
<name>count_up</name></connection>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-25,47.5,-24.5</points>
<connection>
<GID>113</GID>
<name>count_enable</name></connection>
<connection>
<GID>185</GID>
<name>OUT_0</name></connection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>-46.6198,1.65856e-006,35.3604,-89.1089</PageViewport></page 3>
<page 4>
<PageViewport>-46.6198,1.65856e-006,35.3604,-89.1089</PageViewport></page 4>
<page 5>
<PageViewport>-46.6198,1.65856e-006,35.3604,-89.1089</PageViewport></page 5>
<page 6>
<PageViewport>-46.6198,1.65856e-006,35.3604,-89.1089</PageViewport></page 6>
<page 7>
<PageViewport>-46.6198,1.65856e-006,35.3604,-89.1089</PageViewport></page 7>
<page 8>
<PageViewport>-46.6198,1.65856e-006,35.3604,-89.1089</PageViewport></page 8>
<page 9>
<PageViewport>-46.6198,1.65856e-006,35.3604,-89.1089</PageViewport></page 9></circuit>