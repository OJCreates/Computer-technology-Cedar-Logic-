<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-49.4222,20.2,98.4889,-142.17</PageViewport>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>29.5,-9</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_INVERTER</type>
<position>19,-17</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND2</type>
<position>27.5,-26</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>9.5,-25</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Control</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_OR2</type>
<position>45,-17.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>52.5,-17.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>DE_TO</type>
<position>-20.5,-6</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input A</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>-29.5,-6</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>DA_FROM</type>
<position>8,-8</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input A</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_TOGGLE</type>
<position>-29,-19.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>-28.5,-29.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>-19,-19.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Control</lparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>-19,-29.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input B</lparam></gate>
<gate>
<ID>50</ID>
<type>DA_FROM</type>
<position>10.5,-30</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input B</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>9.5,10.5</position>
<gparam>LABEL_TEXT 2-way multiplexer</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>-50.5,-63.5</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>DE_TO</type>
<position>-39.5,-63.5</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input A1</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>-50.5,-74</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>58</ID>
<type>DE_TO</type>
<position>-40,-74</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input B1</lparam></gate>
<gate>
<ID>59</ID>
<type>DE_TO</type>
<position>-39.5,-83</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input A0</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_TOGGLE</type>
<position>-50.5,-83</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>61</ID>
<type>DE_TO</type>
<position>-39,-90.5</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input B0</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>-50,-90.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>-7.5,-59</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input A1</lparam></gate>
<gate>
<ID>65</ID>
<type>DA_FROM</type>
<position>-6,-70.5</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input B1</lparam></gate>
<gate>
<ID>66</ID>
<type>DA_FROM</type>
<position>-6,-77</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input A0</lparam></gate>
<gate>
<ID>67</ID>
<type>DA_FROM</type>
<position>-7,-101.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input B0</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_AND2</type>
<position>35,-58</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>-50.5,-97</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>DE_TO</type>
<position>-38,-96.5</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Control</lparam></gate>
<gate>
<ID>74</ID>
<type>DA_FROM</type>
<position>-7.5,-95</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Control</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_AND2</type>
<position>27.5,-73.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_AND2</type>
<position>28.5,-84.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_AND2</type>
<position>30,-100.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_INVERTER</type>
<position>18.5,-90.5</position>
<input>
<ID>IN_0</ID>31 </input>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>86</ID>
<type>AE_OR2</type>
<position>48.5,-67</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>87</ID>
<type>AE_OR2</type>
<position>47.5,-90</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_TOGGLE</type>
<position>64.5,-66.5</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_TOGGLE</type>
<position>63,-91</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-10,26.5,-10</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>19 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>19,-14,19,-10</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-10 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-25,19,-20</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-25,24.5,-25</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-16.5,37,-9</points>
<intersection>-16.5 1</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-16.5,42,-16.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-9,37,-9</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-26,36,-18.5</points>
<intersection>-26 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-18.5,42,-18.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-26,36,-26</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-17.5,51.5,-17.5</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<connection>
<GID>22</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27.5,-6,-22.5,-6</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-8,26.5,-8</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>26.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>26.5,-8,26.5,-8</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-8 1</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27,-19.5,-21,-19.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-26.5,-29.5,-21,-29.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-30,15.5,-27</points>
<intersection>-30 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,-27,24.5,-27</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-30,15.5,-30</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-48.5,-63.5,-41.5,-63.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-48.5,-74,-42,-74</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-48.5,-83,-41.5,-83</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<connection>
<GID>59</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-48,-90.5,-41,-90.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<connection>
<GID>61</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5.5,-57,32,-57</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>-5.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-5.5,-59,-5.5,-57</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>-57 1</intersection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-97,-44,-96.5</points>
<intersection>-97 2</intersection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-44,-96.5,-40,-96.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>-44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-48.5,-97,-44,-97</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-74.5,10,-70.5</points>
<intersection>-74.5 1</intersection>
<intersection>-70.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-74.5,24.5,-74.5</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4,-70.5,10,-70.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-83.5,11.5,-77</points>
<intersection>-83.5 1</intersection>
<intersection>-77 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-83.5,25.5,-83.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4,-77,11.5,-77</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5,-101.5,27,-101.5</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-99.5,13,-72.5</points>
<intersection>-99.5 2</intersection>
<intersection>-95 3</intersection>
<intersection>-93.5 5</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-72.5,24.5,-72.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-99.5,27,-99.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-5.5,-95,13,-95</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>13,-93.5,18.5,-93.5</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-87.5,18.5,-78</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-78,31,-78</points>
<intersection>18.5 0</intersection>
<intersection>27 3</intersection>
<intersection>31 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>31,-78,31,-59</points>
<intersection>-78 1</intersection>
<intersection>-59 4</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>27,-85.5,27,-78</points>
<intersection>-85.5 5</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>31,-59,32,-59</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>31 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>25.5,-85.5,27,-85.5</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>27 3</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-66,41.5,-58</points>
<intersection>-66 1</intersection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-66,45.5,-66</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-58,41.5,-58</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-89,38,-84.5</points>
<intersection>-89 1</intersection>
<intersection>-84.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-89,44.5,-89</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-84.5,38,-84.5</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-100.5,38.5,-91</points>
<intersection>-100.5 2</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-91,44.5,-91</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-100.5,38.5,-100.5</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-73.5,38,-68</points>
<intersection>-73.5 2</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-68,45.5,-68</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-73.5,38,-73.5</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-67,57,-66.5</points>
<intersection>-67 2</intersection>
<intersection>-66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57,-66.5,62.5,-66.5</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-67,57,-67</points>
<connection>
<GID>86</GID>
<name>OUT</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-91,55.5,-90</points>
<intersection>-91 1</intersection>
<intersection>-90 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-91,61,-91</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-90,55.5,-90</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,62.4,-68.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,62.4,-68.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,62.4,-68.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,62.4,-68.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,62.4,-68.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,62.4,-68.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,62.4,-68.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,62.4,-68.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,62.4,-68.5</PageViewport></page 9></circuit>