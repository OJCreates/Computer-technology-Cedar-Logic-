<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-11.0031,40.0429,141.675,-127.56</PageViewport>
<gate>
<ID>1</ID>
<type>DD_KEYPAD_HEX</type>
<position>42.5,-54.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>2 </output>
<output>
<ID>OUT_3</ID>1 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>2</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>138.5,-55.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>42 </input>
<input>
<ID>IN_2</ID>31 </input>
<input>
<ID>IN_3</ID>32 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>3</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>59.5,-55</position>
<input>
<ID>ENABLE_0</ID>38 </input>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>2 </input>
<input>
<ID>IN_3</ID>1 </input>
<output>
<ID>OUT_0</ID>33 </output>
<output>
<ID>OUT_1</ID>42 </output>
<output>
<ID>OUT_2</ID>31 </output>
<output>
<ID>OUT_3</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_REGISTER4</type>
<position>71,-34.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>42 </input>
<input>
<ID>IN_2</ID>31 </input>
<input>
<ID>IN_3</ID>32 </input>
<output>
<ID>OUT_0</ID>11 </output>
<output>
<ID>OUT_1</ID>9 </output>
<output>
<ID>OUT_2</ID>10 </output>
<output>
<ID>OUT_3</ID>8 </output>
<input>
<ID>clear</ID>7 </input>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>count_enable</ID>6 </input>
<input>
<ID>count_up</ID>5 </input>
<input>
<ID>load</ID>14 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>5</ID>
<type>FF_GND</type>
<position>72,-28.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>FF_GND</type>
<position>71,-27</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>FF_GND</type>
<position>72,-39.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>77.5,-34</position>
<input>
<ID>ENABLE_0</ID>39 </input>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>9 </input>
<input>
<ID>IN_2</ID>10 </input>
<input>
<ID>IN_3</ID>8 </input>
<output>
<ID>OUT_0</ID>33 </output>
<output>
<ID>OUT_1</ID>42 </output>
<output>
<ID>OUT_2</ID>31 </output>
<output>
<ID>OUT_3</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>9</ID>
<type>DA_FROM</type>
<position>70,-40.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>10</ID>
<type>DE_TO</type>
<position>47.5,-67.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>41.5,-67.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>BA_DECODER_2x4</type>
<position>55,-22</position>
<input>
<ID>ENABLE</ID>36 </input>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT_1</ID>14 </output>
<output>
<ID>OUT_2</ID>34 </output>
<output>
<ID>OUT_3</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_REGISTER4</type>
<position>93,-34.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>42 </input>
<input>
<ID>IN_2</ID>31 </input>
<input>
<ID>IN_3</ID>32 </input>
<output>
<ID>OUT_0</ID>21 </output>
<output>
<ID>OUT_1</ID>19 </output>
<output>
<ID>OUT_2</ID>20 </output>
<output>
<ID>OUT_3</ID>18 </output>
<input>
<ID>clear</ID>17 </input>
<input>
<ID>clock</ID>22 </input>
<input>
<ID>count_enable</ID>16 </input>
<input>
<ID>count_up</ID>15 </input>
<input>
<ID>load</ID>34 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>14</ID>
<type>FF_GND</type>
<position>94,-28.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>FF_GND</type>
<position>93,-27</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>FF_GND</type>
<position>94,-39.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>99.5,-34</position>
<input>
<ID>ENABLE_0</ID>40 </input>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>19 </input>
<input>
<ID>IN_2</ID>20 </input>
<input>
<ID>IN_3</ID>18 </input>
<output>
<ID>OUT_0</ID>33 </output>
<output>
<ID>OUT_1</ID>42 </output>
<output>
<ID>OUT_2</ID>31 </output>
<output>
<ID>OUT_3</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>92,-40.5</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_REGISTER4</type>
<position>120.5,-34.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>42 </input>
<input>
<ID>IN_2</ID>31 </input>
<input>
<ID>IN_3</ID>32 </input>
<output>
<ID>OUT_0</ID>29 </output>
<output>
<ID>OUT_1</ID>27 </output>
<output>
<ID>OUT_2</ID>28 </output>
<output>
<ID>OUT_3</ID>26 </output>
<input>
<ID>clear</ID>25 </input>
<input>
<ID>clock</ID>30 </input>
<input>
<ID>count_enable</ID>24 </input>
<input>
<ID>count_up</ID>23 </input>
<input>
<ID>load</ID>35 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 8</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>20</ID>
<type>FF_GND</type>
<position>121.5,-28.5</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>21</ID>
<type>FF_GND</type>
<position>120.5,-27</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>FF_GND</type>
<position>121.5,-39.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>23</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>127,-34</position>
<input>
<ID>ENABLE_0</ID>41 </input>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>27 </input>
<input>
<ID>IN_2</ID>28 </input>
<input>
<ID>IN_3</ID>26 </input>
<output>
<ID>OUT_0</ID>33 </output>
<output>
<ID>OUT_1</ID>42 </output>
<output>
<ID>OUT_2</ID>31 </output>
<output>
<ID>OUT_3</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>119.5,-40.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>25</ID>
<type>BA_DECODER_2x4</type>
<position>54.5,-15.5</position>
<input>
<ID>ENABLE</ID>37 </input>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT_0</ID>38 </output>
<output>
<ID>OUT_1</ID>39 </output>
<output>
<ID>OUT_2</ID>40 </output>
<output>
<ID>OUT_3</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>EE_VDD</type>
<position>50.5,-14</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>27</ID>
<type>EE_VDD</type>
<position>50,-21.5</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AE_REGISTER8</type>
<position>32,-22</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>74 </input>
<input>
<ID>IN_2</ID>75 </input>
<input>
<ID>IN_3</ID>76 </input>
<input>
<ID>IN_4</ID>77 </input>
<input>
<ID>IN_5</ID>78 </input>
<input>
<ID>IN_6</ID>79 </input>
<input>
<ID>IN_7</ID>80 </input>
<output>
<ID>OUT_0</ID>59 </output>
<output>
<ID>OUT_1</ID>58 </output>
<output>
<ID>OUT_2</ID>57 </output>
<output>
<ID>OUT_3</ID>56 </output>
<output>
<ID>OUT_4</ID>46 </output>
<output>
<ID>OUT_5</ID>45 </output>
<output>
<ID>OUT_6</ID>44 </output>
<output>
<ID>OUT_7</ID>43 </output>
<input>
<ID>clear</ID>48 </input>
<input>
<ID>clock</ID>47 </input>
<input>
<ID>count_enable</ID>49 </input>
<input>
<ID>count_up</ID>49 </input>
<input>
<ID>load</ID>50 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 180</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>29</ID>
<type>DA_FROM</type>
<position>31,-32</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Clock</lparam></gate>
<gate>
<ID>30</ID>
<type>FF_GND</type>
<position>33,-28</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>FF_GND</type>
<position>33,-13.5</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>EE_VDD</type>
<position>31,-13</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>33</ID>
<type>BA_ROM_4x4</type>
<position>6.5,-15</position>
<input>
<ID>ADDRESS_0</ID>63 </input>
<input>
<ID>ADDRESS_1</ID>62 </input>
<input>
<ID>ADDRESS_2</ID>61 </input>
<input>
<ID>ADDRESS_3</ID>60 </input>
<output>
<ID>DATA_OUT_0</ID>77 </output>
<output>
<ID>DATA_OUT_1</ID>78 </output>
<output>
<ID>DATA_OUT_2</ID>79 </output>
<output>
<ID>DATA_OUT_3</ID>80 </output>
<input>
<ID>ENABLE_0</ID>55 </input>
<gparam>angle 90</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:0 1</lparam>
<lparam>Address:1 6</lparam>
<lparam>Address:2 1</lparam>
<lparam>Address:3 11</lparam></gate>
<gate>
<ID>34</ID>
<type>EE_VDD</type>
<position>7,-8</position>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>35</ID>
<type>DE_TO</type>
<position>47,-26.5</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>36</ID>
<type>DE_TO</type>
<position>47,-29.5</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>37</ID>
<type>DE_TO</type>
<position>47,-33</position>
<input>
<ID>IN_0</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>38</ID>
<type>DE_TO</type>
<position>47,-36</position>
<input>
<ID>IN_0</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>39</ID>
<type>DA_FROM</type>
<position>3,-24.5</position>
<input>
<ID>IN_0</ID>60 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>40</ID>
<type>DA_FROM</type>
<position>5.5,-24.5</position>
<input>
<ID>IN_0</ID>61 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>41</ID>
<type>DA_FROM</type>
<position>8,-24.5</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>10.5,-24.5</position>
<input>
<ID>IN_0</ID>63 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>43</ID>
<type>BA_ROM_4x4</type>
<position>6,-33.5</position>
<input>
<ID>ADDRESS_0</ID>68 </input>
<input>
<ID>ADDRESS_1</ID>67 </input>
<input>
<ID>ADDRESS_2</ID>66 </input>
<input>
<ID>ADDRESS_3</ID>65 </input>
<output>
<ID>DATA_OUT_0</ID>73 </output>
<output>
<ID>DATA_OUT_1</ID>74 </output>
<output>
<ID>DATA_OUT_2</ID>75 </output>
<output>
<ID>DATA_OUT_3</ID>76 </output>
<input>
<ID>ENABLE_0</ID>64 </input>
<gparam>angle 90</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:0 1</lparam>
<lparam>Address:1 2</lparam>
<lparam>Address:2 3</lparam>
<lparam>Address:3 4</lparam></gate>
<gate>
<ID>44</ID>
<type>EE_VDD</type>
<position>6.5,-27.5</position>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>45</ID>
<type>DA_FROM</type>
<position>3,-57</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>46</ID>
<type>DA_FROM</type>
<position>5.5,-57</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>47</ID>
<type>DA_FROM</type>
<position>8,-57</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>48</ID>
<type>DA_FROM</type>
<position>10.5,-57</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-53.5,52.5,-51.5</points>
<intersection>-53.5 5</intersection>
<intersection>-51.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>47.5,-51.5,52.5,-51.5</points>
<connection>
<GID>1</GID>
<name>OUT_3</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>52.5,-53.5,57.5,-53.5</points>
<connection>
<GID>3</GID>
<name>IN_3</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-54.5,52.5,-53.5</points>
<intersection>-54.5 4</intersection>
<intersection>-53.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47.5,-53.5,52.5,-53.5</points>
<connection>
<GID>1</GID>
<name>OUT_2</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52.5,-54.5,57.5,-54.5</points>
<connection>
<GID>3</GID>
<name>IN_2</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>47.5,-55.5,57.5,-55.5</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<connection>
<GID>1</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-57.5,52.5,-56.5</points>
<intersection>-57.5 3</intersection>
<intersection>-56.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47.5,-57.5,52.5,-57.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52.5,-56.5,57.5,-56.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>72,-29.5,72,-29.5</points>
<connection>
<GID>4</GID>
<name>count_up</name></connection>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-29.5,71,-28</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>4</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>72,-38.5,72,-38.5</points>
<connection>
<GID>4</GID>
<name>clear</name></connection>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>75,-32.5,75.5,-32.5</points>
<connection>
<GID>8</GID>
<name>IN_3</name></connection>
<connection>
<GID>4</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>75,-34.5,75.5,-34.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<connection>
<GID>4</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>75,-33.5,75.5,-33.5</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<connection>
<GID>4</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>75,-35.5,75.5,-35.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>70,-38.5,70,-38.5</points>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<connection>
<GID>9</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43.5,-67.5,45.5,-67.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-29.5,70,-22.5</points>
<connection>
<GID>4</GID>
<name>load</name></connection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-22.5,70,-22.5</points>
<connection>
<GID>12</GID>
<name>OUT_1</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>94,-29.5,94,-29.5</points>
<connection>
<GID>13</GID>
<name>count_up</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-29.5,93,-28</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<connection>
<GID>13</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>94,-38.5,94,-38.5</points>
<connection>
<GID>13</GID>
<name>clear</name></connection>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97,-32.5,97.5,-32.5</points>
<connection>
<GID>17</GID>
<name>IN_3</name></connection>
<connection>
<GID>13</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97,-34.5,97.5,-34.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<connection>
<GID>13</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97,-33.5,97.5,-33.5</points>
<connection>
<GID>17</GID>
<name>IN_2</name></connection>
<connection>
<GID>13</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97,-35.5,97.5,-35.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>92,-38.5,92,-38.5</points>
<connection>
<GID>13</GID>
<name>clock</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-29.5,121.5,-29.5</points>
<connection>
<GID>19</GID>
<name>count_up</name></connection>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120.5,-29.5,120.5,-28</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<connection>
<GID>19</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-38.5,121.5,-38.5</points>
<connection>
<GID>19</GID>
<name>clear</name></connection>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124.5,-32.5,125,-32.5</points>
<connection>
<GID>23</GID>
<name>IN_3</name></connection>
<connection>
<GID>19</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124.5,-34.5,125,-34.5</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<connection>
<GID>19</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124.5,-33.5,125,-33.5</points>
<connection>
<GID>23</GID>
<name>IN_2</name></connection>
<connection>
<GID>19</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124.5,-35.5,125,-35.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>119.5,-38.5,119.5,-38.5</points>
<connection>
<GID>19</GID>
<name>clock</name></connection>
<connection>
<GID>24</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61.5,-54.5,135.5,-54.5</points>
<connection>
<GID>3</GID>
<name>OUT_2</name></connection>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>65 8</intersection>
<intersection>81.5 12</intersection>
<intersection>87 13</intersection>
<intersection>104.5 20</intersection>
<intersection>114.5 21</intersection>
<intersection>131 19</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>65,-54.5,65,-33.5</points>
<intersection>-54.5 1</intersection>
<intersection>-33.5 25</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>81.5,-54.5,81.5,-33.5</points>
<intersection>-54.5 1</intersection>
<intersection>-33.5 16</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>87,-54.5,87,-33.5</points>
<intersection>-54.5 1</intersection>
<intersection>-33.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>87,-33.5,89,-33.5</points>
<connection>
<GID>13</GID>
<name>IN_2</name></connection>
<intersection>87 13</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>79.5,-33.5,81.5,-33.5</points>
<connection>
<GID>8</GID>
<name>OUT_2</name></connection>
<intersection>81.5 12</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>131,-54.5,131,-33.5</points>
<intersection>-54.5 1</intersection>
<intersection>-33.5 24</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>104.5,-54.5,104.5,-33.5</points>
<intersection>-54.5 1</intersection>
<intersection>-33.5 22</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>114.5,-54.5,114.5,-33.5</points>
<intersection>-54.5 1</intersection>
<intersection>-33.5 23</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>101.5,-33.5,104.5,-33.5</points>
<connection>
<GID>17</GID>
<name>OUT_2</name></connection>
<intersection>104.5 20</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>114.5,-33.5,116.5,-33.5</points>
<connection>
<GID>19</GID>
<name>IN_2</name></connection>
<intersection>114.5 21</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>129,-33.5,131,-33.5</points>
<connection>
<GID>23</GID>
<name>OUT_2</name></connection>
<intersection>131 19</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>65,-33.5,67,-33.5</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<intersection>65 8</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61.5,-53.5,135.5,-53.5</points>
<connection>
<GID>3</GID>
<name>OUT_3</name></connection>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>63.5 9</intersection>
<intersection>82 13</intersection>
<intersection>85.5 14</intersection>
<intersection>105.5 23</intersection>
<intersection>113.5 24</intersection>
<intersection>132.5 22</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>63.5,-53.5,63.5,-32.5</points>
<intersection>-53.5 1</intersection>
<intersection>-32.5 29</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>82,-53.5,82,-32.5</points>
<intersection>-53.5 1</intersection>
<intersection>-32.5 28</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>85.5,-53.5,85.5,-32.5</points>
<intersection>-53.5 1</intersection>
<intersection>-32.5 20</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>85.5,-32.5,89,-32.5</points>
<connection>
<GID>13</GID>
<name>IN_3</name></connection>
<intersection>85.5 14</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>132.5,-53.5,132.5,-32.5</points>
<intersection>-53.5 1</intersection>
<intersection>-32.5 27</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>105.5,-53.5,105.5,-32.5</points>
<intersection>-53.5 1</intersection>
<intersection>-32.5 25</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>113.5,-53.5,113.5,-32.5</points>
<intersection>-53.5 1</intersection>
<intersection>-32.5 26</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>101.5,-32.5,105.5,-32.5</points>
<connection>
<GID>17</GID>
<name>OUT_3</name></connection>
<intersection>105.5 23</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>113.5,-32.5,116.5,-32.5</points>
<connection>
<GID>19</GID>
<name>IN_3</name></connection>
<intersection>113.5 24</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>129,-32.5,132.5,-32.5</points>
<connection>
<GID>23</GID>
<name>OUT_3</name></connection>
<intersection>132.5 22</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>79.5,-32.5,82,-32.5</points>
<connection>
<GID>8</GID>
<name>OUT_3</name></connection>
<intersection>82 13</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>63.5,-32.5,67,-32.5</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<intersection>63.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61.5,-56.5,135.5,-56.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>67 4</intersection>
<intersection>79.5 6</intersection>
<intersection>89 10</intersection>
<intersection>101.5 9</intersection>
<intersection>116.5 14</intersection>
<intersection>129 13</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>67,-56.5,67,-35.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>79.5,-56.5,79.5,-35.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>101.5,-56.5,101.5,-35.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>89,-56.5,89,-35.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>129,-56.5,129,-35.5</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>116.5,-56.5,116.5,-35.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-56.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-29.5,92,-21.5</points>
<connection>
<GID>13</GID>
<name>load</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-21.5,92,-21.5</points>
<connection>
<GID>12</GID>
<name>OUT_2</name></connection>
<intersection>92 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-29.5,119.5,-20.5</points>
<connection>
<GID>19</GID>
<name>load</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-20.5,119.5,-20.5</points>
<connection>
<GID>12</GID>
<name>OUT_3</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-21.5,52,-20.5</points>
<connection>
<GID>12</GID>
<name>ENABLE</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-21.5,52,-21.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>51.5,-14,51.5,-14</points>
<connection>
<GID>25</GID>
<name>ENABLE</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-52,59.5,-17</points>
<connection>
<GID>3</GID>
<name>ENABLE_0</name></connection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-17,59.5,-17</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-31,77.5,-16</points>
<connection>
<GID>8</GID>
<name>ENABLE_0</name></connection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-16,77.5,-16</points>
<connection>
<GID>25</GID>
<name>OUT_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-31,99.5,-15</points>
<connection>
<GID>17</GID>
<name>ENABLE_0</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-15,99.5,-15</points>
<connection>
<GID>25</GID>
<name>OUT_2</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-31,127,-14</points>
<connection>
<GID>23</GID>
<name>ENABLE_0</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-14,127,-14</points>
<connection>
<GID>25</GID>
<name>OUT_3</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61.5,-55.5,135.5,-55.5</points>
<connection>
<GID>3</GID>
<name>OUT_1</name></connection>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>66 7</intersection>
<intersection>80.5 12</intersection>
<intersection>88 13</intersection>
<intersection>103 20</intersection>
<intersection>115.5 21</intersection>
<intersection>130 19</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>66,-55.5,66,-34.5</points>
<intersection>-55.5 1</intersection>
<intersection>-34.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>66,-34.5,67,-34.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>66 7</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>80.5,-55.5,80.5,-34.5</points>
<intersection>-55.5 1</intersection>
<intersection>-34.5 16</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>88,-55.5,88,-34.5</points>
<intersection>-55.5 1</intersection>
<intersection>-34.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>88,-34.5,89,-34.5</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>88 13</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>79.5,-34.5,80.5,-34.5</points>
<connection>
<GID>8</GID>
<name>OUT_1</name></connection>
<intersection>80.5 12</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>130,-55.5,130,-34.5</points>
<intersection>-55.5 1</intersection>
<intersection>-34.5 24</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>103,-55.5,103,-34.5</points>
<intersection>-55.5 1</intersection>
<intersection>-34.5 22</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>115.5,-55.5,115.5,-34.5</points>
<intersection>-55.5 1</intersection>
<intersection>-34.5 23</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>101.5,-34.5,103,-34.5</points>
<connection>
<GID>17</GID>
<name>OUT_1</name></connection>
<intersection>103 20</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>115.5,-34.5,116.5,-34.5</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>115.5 21</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>129,-34.5,130,-34.5</points>
<connection>
<GID>23</GID>
<name>OUT_1</name></connection>
<intersection>130 19</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-18,43.5,-16</points>
<intersection>-18 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-16,51.5,-16</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36,-18,43.5,-18</points>
<connection>
<GID>28</GID>
<name>OUT_7</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-19,44.5,-17</points>
<intersection>-19 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-17,51.5,-17</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36,-19,44.5,-19</points>
<connection>
<GID>28</GID>
<name>OUT_6</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-22.5,45,-20</points>
<intersection>-22.5 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-22.5,52,-22.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36,-20,45,-20</points>
<connection>
<GID>28</GID>
<name>OUT_5</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-23.5,44,-21</points>
<intersection>-23.5 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-23.5,52,-23.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36,-21,44,-21</points>
<connection>
<GID>28</GID>
<name>OUT_4</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-30,31,-27</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-27,33,-27</points>
<connection>
<GID>28</GID>
<name>clear</name></connection>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-16,33,-14.5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<connection>
<GID>28</GID>
<name>count_up</name></connection>
<intersection>-16 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>32,-16,33,-16</points>
<connection>
<GID>28</GID>
<name>count_enable</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-16,31,-14</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<connection>
<GID>28</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-10,7,-9</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<connection>
<GID>33</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-26.5,43,-22</points>
<intersection>-26.5 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-22,43,-22</points>
<connection>
<GID>28</GID>
<name>OUT_3</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-26.5,45,-26.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-29.5,41.5,-23</points>
<intersection>-29.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-23,41.5,-23</points>
<connection>
<GID>28</GID>
<name>OUT_2</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-29.5,45,-29.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-33,40.5,-24</points>
<intersection>-33 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-24,40.5,-24</points>
<connection>
<GID>28</GID>
<name>OUT_1</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-33,45,-33</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-36,39,-25</points>
<intersection>-36 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-36,45,-36</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36,-25,39,-25</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-21.5,5,-20</points>
<connection>
<GID>33</GID>
<name>ADDRESS_3</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>3,-22.5,3,-21.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>3,-21.5,5,-21.5</points>
<intersection>3 1</intersection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-21.5,6,-20</points>
<connection>
<GID>33</GID>
<name>ADDRESS_2</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>5.5,-22.5,5.5,-21.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>5.5,-21.5,6,-21.5</points>
<intersection>5.5 1</intersection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-21.5,7,-20</points>
<connection>
<GID>33</GID>
<name>ADDRESS_1</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>8,-22.5,8,-21.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>7,-21.5,8,-21.5</points>
<intersection>7 0</intersection>
<intersection>8 1</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-21,8,-20</points>
<connection>
<GID>33</GID>
<name>ADDRESS_0</name></connection>
<intersection>-21 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>10.5,-22.5,10.5,-21</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>8,-21,10.5,-21</points>
<intersection>8 0</intersection>
<intersection>10.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-28.5,6.5,-28.5</points>
<connection>
<GID>43</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-51,4.5,-38.5</points>
<connection>
<GID>43</GID>
<name>ADDRESS_3</name></connection>
<intersection>-51 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>3,-55,3,-51</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>3,-51,4.5,-51</points>
<intersection>3 1</intersection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-55,5.5,-38.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<connection>
<GID>43</GID>
<name>ADDRESS_2</name></connection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-48,6.5,-38.5</points>
<connection>
<GID>43</GID>
<name>ADDRESS_1</name></connection>
<intersection>-48 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>8,-55,8,-48</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-48,8,-48</points>
<intersection>6.5 0</intersection>
<intersection>8 1</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-46,7.5,-38.5</points>
<connection>
<GID>43</GID>
<name>ADDRESS_0</name></connection>
<intersection>-46 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>10.5,-55,10.5,-46</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-46,10.5,-46</points>
<intersection>7.5 0</intersection>
<intersection>10.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-32,17,-25</points>
<intersection>-32 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-25,28,-25</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-32,17,-32</points>
<connection>
<GID>43</GID>
<name>DATA_OUT_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-33,19.5,-24</points>
<intersection>-33 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-24,28,-24</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-33,19.5,-33</points>
<connection>
<GID>43</GID>
<name>DATA_OUT_1</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-34,21.5,-23</points>
<intersection>-34 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-23,28,-23</points>
<connection>
<GID>28</GID>
<name>IN_2</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-34,21.5,-34</points>
<connection>
<GID>43</GID>
<name>DATA_OUT_2</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-35,23.5,-22</points>
<intersection>-35 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-22,28,-22</points>
<connection>
<GID>28</GID>
<name>IN_3</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-35,23.5,-35</points>
<connection>
<GID>43</GID>
<name>DATA_OUT_3</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-21,23.5,-13.5</points>
<intersection>-21 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-21,28,-21</points>
<connection>
<GID>28</GID>
<name>IN_4</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-13.5,23.5,-13.5</points>
<connection>
<GID>33</GID>
<name>DATA_OUT_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-20,21.5,-14.5</points>
<intersection>-20 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-20,28,-20</points>
<connection>
<GID>28</GID>
<name>IN_5</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-14.5,21.5,-14.5</points>
<connection>
<GID>33</GID>
<name>DATA_OUT_1</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-19,19.5,-15.5</points>
<intersection>-19 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-19,28,-19</points>
<connection>
<GID>28</GID>
<name>IN_6</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-15.5,19.5,-15.5</points>
<connection>
<GID>33</GID>
<name>DATA_OUT_2</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-18,16.5,-16.5</points>
<intersection>-18 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-18,28,-18</points>
<connection>
<GID>28</GID>
<name>IN_7</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-16.5,16.5,-16.5</points>
<connection>
<GID>33</GID>
<name>DATA_OUT_3</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,189.465,482.538,-340.244</PageViewport></page 1>
<page 2>
<PageViewport>0,189.465,482.538,-340.244</PageViewport></page 2>
<page 3>
<PageViewport>0,189.465,482.538,-340.244</PageViewport></page 3>
<page 4>
<PageViewport>0,189.465,482.538,-340.244</PageViewport></page 4>
<page 5>
<PageViewport>0,189.465,482.538,-340.244</PageViewport></page 5>
<page 6>
<PageViewport>0,189.465,482.538,-340.244</PageViewport></page 6>
<page 7>
<PageViewport>0,189.465,482.538,-340.244</PageViewport></page 7>
<page 8>
<PageViewport>0,189.465,482.538,-340.244</PageViewport></page 8>
<page 9>
<PageViewport>0,189.465,482.538,-340.244</PageViewport></page 9></circuit>