<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>14.4556,14.4296,159.522,-145.57</PageViewport>
<gate>
<ID>2</ID>
<type>DD_KEYPAD_HEX</type>
<position>23.5,-42.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<output>
<ID>OUT_1</ID>9 </output>
<output>
<ID>OUT_2</ID>7 </output>
<output>
<ID>OUT_3</ID>6 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>3</ID>
<type>DD_KEYPAD_HEX</type>
<position>63.5,-13.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<output>
<ID>OUT_1</ID>27 </output>
<output>
<ID>OUT_2</ID>26 </output>
<output>
<ID>OUT_3</ID>25 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 13</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_FULLADDER_4BIT</type>
<position>42,-61</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>12 </input>
<input>
<ID>IN_2</ID>11 </input>
<input>
<ID>IN_3</ID>10 </input>
<input>
<ID>IN_B_0</ID>24 </input>
<input>
<ID>IN_B_1</ID>23 </input>
<input>
<ID>IN_B_2</ID>22 </input>
<input>
<ID>IN_B_3</ID>21 </input>
<output>
<ID>OUT_0</ID>16 </output>
<output>
<ID>OUT_1</ID>17 </output>
<output>
<ID>OUT_2</ID>18 </output>
<output>
<ID>OUT_3</ID>19 </output>
<input>
<ID>carry_in</ID>33 </input>
<output>
<ID>carry_out</ID>14 </output>
<output>
<ID>overflow</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>9</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>38.5,-43</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>6 </input>
<output>
<ID>OUT_0</ID>13 </output>
<output>
<ID>OUT_1</ID>12 </output>
<output>
<ID>OUT_2</ID>11 </output>
<output>
<ID>OUT_3</ID>10 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>11</ID>
<type>GA_LED</type>
<position>24,-57.5</position>
<input>
<ID>N_in1</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>24,-62.5</position>
<input>
<ID>N_in1</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>32,-74</position>
<input>
<ID>N_in1</ID>19 </input>
<input>
<ID>N_in2</ID>20 </input>
<input>
<ID>N_in3</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>47.5,-71.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>17 </input>
<input>
<ID>IN_2</ID>18 </input>
<input>
<ID>IN_3</ID>19 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>18</ID>
<type>AI_XOR2</type>
<position>65.5,-41</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AI_XOR2</type>
<position>75.5,-41</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AI_XOR2</type>
<position>87,-41</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>AI_XOR2</type>
<position>98,-41</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>81.5,-14</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>27 </input>
<input>
<ID>IN_2</ID>26 </input>
<input>
<ID>IN_3</ID>25 </input>
<output>
<ID>OUT_0</ID>32 </output>
<output>
<ID>OUT_1</ID>31 </output>
<output>
<ID>OUT_2</ID>30 </output>
<output>
<ID>OUT_3</ID>29 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 13</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>23</ID>
<type>AE_FULLADDER_4BIT</type>
<position>147,-61</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>37 </input>
<input>
<ID>IN_3</ID>36 </input>
<input>
<ID>IN_B_0</ID>51 </input>
<input>
<ID>IN_B_1</ID>50 </input>
<input>
<ID>IN_B_2</ID>49 </input>
<input>
<ID>IN_B_3</ID>48 </input>
<output>
<ID>OUT_0</ID>47 </output>
<output>
<ID>OUT_1</ID>46 </output>
<output>
<ID>OUT_2</ID>45 </output>
<output>
<ID>OUT_3</ID>44 </output>
<input>
<ID>carry_in</ID>53 </input>
<output>
<ID>carry_out</ID>33 </output>
<output>
<ID>overflow</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>25</ID>
<type>GA_LED</type>
<position>132.5,-64.5</position>
<input>
<ID>N_in1</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>143.5,-44</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>42 </input>
<input>
<ID>IN_2</ID>41 </input>
<input>
<ID>IN_3</ID>40 </input>
<output>
<ID>OUT_0</ID>39 </output>
<output>
<ID>OUT_1</ID>38 </output>
<output>
<ID>OUT_2</ID>37 </output>
<output>
<ID>OUT_3</ID>36 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>28</ID>
<type>DD_KEYPAD_HEX</type>
<position>128,-43</position>
<output>
<ID>OUT_0</ID>43 </output>
<output>
<ID>OUT_1</ID>42 </output>
<output>
<ID>OUT_2</ID>41 </output>
<output>
<ID>OUT_3</ID>40 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 7</lparam></gate>
<gate>
<ID>30</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>153.5,-73</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>46 </input>
<input>
<ID>IN_2</ID>45 </input>
<input>
<ID>IN_3</ID>44 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>31</ID>
<type>AI_XOR2</type>
<position>160,-42</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AI_XOR2</type>
<position>170,-42</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>AI_XOR2</type>
<position>180,-42</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>AI_XOR2</type>
<position>189,-42</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>202,-34.5</position>
<input>
<ID>IN_0</ID>53 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Add/Sub</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>151.5,-92.5</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>165.5,-92</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Add/Sub</lparam></gate>
<gate>
<ID>41</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>169.5,-17.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>61 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>58 </input>
<output>
<ID>OUT_0</ID>57 </output>
<output>
<ID>OUT_1</ID>56 </output>
<output>
<ID>OUT_2</ID>55 </output>
<output>
<ID>OUT_3</ID>54 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>42</ID>
<type>DD_KEYPAD_HEX</type>
<position>140,-17</position>
<output>
<ID>OUT_0</ID>60 </output>
<output>
<ID>OUT_1</ID>61 </output>
<output>
<ID>OUT_2</ID>59 </output>
<output>
<ID>OUT_3</ID>58 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 9</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>133.5,-68.5</position>
<gparam>LABEL_TEXT Overflow</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>32.5,-78</position>
<gparam>LABEL_TEXT Negative</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>15,-56.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-41,32,-39.5</points>
<intersection>-41 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-39.5,32,-39.5</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-41,35.5,-41</points>
<connection>
<GID>9</GID>
<name>IN_3</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-42,32,-41.5</points>
<intersection>-42 2</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-41.5,32,-41.5</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-42,35.5,-42</points>
<connection>
<GID>9</GID>
<name>IN_2</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-45.5,32,-44</points>
<intersection>-45.5 1</intersection>
<intersection>-44 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-45.5,32,-45.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-44,35.5,-44</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-43.5,32,-43</points>
<intersection>-43.5 1</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-43.5,32,-43.5</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-43,35.5,-43</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-57,37,-47</points>
<connection>
<GID>7</GID>
<name>IN_3</name></connection>
<connection>
<GID>9</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-57,38,-47</points>
<connection>
<GID>7</GID>
<name>IN_2</name></connection>
<connection>
<GID>9</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-57,39,-47</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<connection>
<GID>9</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-57,40,-47</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-60,29.5,-57.5</points>
<intersection>-60 2</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-57.5,29.5,-57.5</points>
<connection>
<GID>11</GID>
<name>N_in1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-60,34,-60</points>
<connection>
<GID>7</GID>
<name>carry_out</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-62.5,34,-62.5</points>
<connection>
<GID>12</GID>
<name>N_in1</name></connection>
<intersection>34 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34,-62.5,34,-62</points>
<connection>
<GID>7</GID>
<name>overflow</name></connection>
<intersection>-62.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-72.5,43.5,-65</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-72.5,44.5,-72.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-71.5,42.5,-65</points>
<connection>
<GID>7</GID>
<name>OUT_1</name></connection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-71.5,44.5,-71.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-70.5,41.5,-65</points>
<connection>
<GID>7</GID>
<name>OUT_2</name></connection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-70.5,44.5,-70.5</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-74,40.5,-65</points>
<connection>
<GID>7</GID>
<name>OUT_3</name></connection>
<intersection>-74 2</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-69.5,44.5,-69.5</points>
<connection>
<GID>16</GID>
<name>IN_3</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-74,40.5,-74</points>
<connection>
<GID>14</GID>
<name>N_in1</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-75,31.5,-73</points>
<intersection>-75 4</intersection>
<intersection>-73 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-73,32,-73</points>
<connection>
<GID>14</GID>
<name>N_in3</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>31.5,-75,32,-75</points>
<connection>
<GID>14</GID>
<name>N_in2</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-50.5,65.5,-44</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>-50.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>44,-57,44,-50.5</points>
<connection>
<GID>7</GID>
<name>IN_B_3</name></connection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>44,-50.5,65.5,-50.5</points>
<intersection>44 1</intersection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-52,75.5,-44</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>-52 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>45,-57,45,-52</points>
<connection>
<GID>7</GID>
<name>IN_B_2</name></connection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45,-52,75.5,-52</points>
<intersection>45 1</intersection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-53.5,87,-44</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>46,-57,46,-53.5</points>
<connection>
<GID>7</GID>
<name>IN_B_1</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>46,-53.5,87,-53.5</points>
<intersection>46 1</intersection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-54.5,98,-44</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<intersection>-54.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>47,-57,47,-54.5</points>
<connection>
<GID>7</GID>
<name>IN_B_0</name></connection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47,-54.5,98,-54.5</points>
<intersection>47 1</intersection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-12,73.5,-10.5</points>
<intersection>-12 1</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-12,78.5,-12</points>
<connection>
<GID>22</GID>
<name>IN_3</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68.5,-10.5,73.5,-10.5</points>
<connection>
<GID>3</GID>
<name>OUT_3</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68.5,-12.5,78.5,-12.5</points>
<connection>
<GID>3</GID>
<name>OUT_2</name></connection>
<intersection>78.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-13,78.5,-12.5</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-14.5,73.5,-14</points>
<intersection>-14.5 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-14.5,73.5,-14.5</points>
<connection>
<GID>3</GID>
<name>OUT_1</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-14,78.5,-14</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-16.5,73.5,-15</points>
<intersection>-16.5 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-16.5,73.5,-16.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-15,78.5,-15</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-38,64.5,-28</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>-28 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>80,-28,80,-18</points>
<connection>
<GID>22</GID>
<name>OUT_3</name></connection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-28,80,-28</points>
<intersection>64.5 0</intersection>
<intersection>80 1</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-38,74.5,-30.5</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>-30.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>81,-30.5,81,-18</points>
<connection>
<GID>22</GID>
<name>OUT_2</name></connection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-30.5,81,-30.5</points>
<intersection>74.5 0</intersection>
<intersection>81 1</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-38,86,-28</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>-28 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>82,-28,82,-18</points>
<connection>
<GID>22</GID>
<name>OUT_1</name></connection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>82,-28,86,-28</points>
<intersection>82 1</intersection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-38,97,-28</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>-28 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>83,-28,83,-18</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>83,-28,97,-28</points>
<intersection>83 1</intersection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-60,139,-60</points>
<connection>
<GID>7</GID>
<name>carry_in</name></connection>
<connection>
<GID>23</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-64.5,136,-62</points>
<intersection>-64.5 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136,-62,139,-62</points>
<connection>
<GID>23</GID>
<name>overflow</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>133.5,-64.5,136,-64.5</points>
<connection>
<GID>25</GID>
<name>N_in1</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-57,142,-48</points>
<connection>
<GID>23</GID>
<name>IN_3</name></connection>
<connection>
<GID>26</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-57,143,-48</points>
<connection>
<GID>23</GID>
<name>IN_2</name></connection>
<connection>
<GID>26</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-57,144,-48</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<connection>
<GID>26</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-57,145,-48</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-40.5,140.5,-40.5</points>
<intersection>133 4</intersection>
<intersection>140.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>140.5,-42,140.5,-40.5</points>
<connection>
<GID>26</GID>
<name>IN_3</name></connection>
<intersection>-40.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>133,-40.5,133,-40</points>
<intersection>-40.5 1</intersection>
<intersection>-40 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>133,-40,133,-40</points>
<connection>
<GID>28</GID>
<name>OUT_3</name></connection>
<intersection>133 4</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-43,140.5,-43</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>133 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>133,-43,133,-42</points>
<intersection>-43 1</intersection>
<intersection>-42 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>133,-42,133,-42</points>
<connection>
<GID>28</GID>
<name>OUT_2</name></connection>
<intersection>133 7</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-44,140.5,-44</points>
<connection>
<GID>28</GID>
<name>OUT_1</name></connection>
<intersection>140.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>140.5,-44,140.5,-44</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-45,140.5,-45</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>133 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>133,-46,133,-45</points>
<intersection>-46 6</intersection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>133,-46,133,-46</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>133 5</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-71,145.5,-65</points>
<connection>
<GID>23</GID>
<name>OUT_3</name></connection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,-71,150.5,-71</points>
<connection>
<GID>30</GID>
<name>IN_3</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-72,146.5,-65</points>
<connection>
<GID>23</GID>
<name>OUT_2</name></connection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>146.5,-72,150.5,-72</points>
<connection>
<GID>30</GID>
<name>IN_2</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,-73,147.5,-65</points>
<connection>
<GID>23</GID>
<name>OUT_1</name></connection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147.5,-73,150.5,-73</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-74,148.5,-65</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148.5,-74,150.5,-74</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>148.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-51,160,-45</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>-51 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>149,-57,149,-51</points>
<connection>
<GID>23</GID>
<name>IN_B_3</name></connection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>149,-51,160,-51</points>
<intersection>149 1</intersection>
<intersection>160 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-51,170,-45</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<intersection>-51 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>150,-57,150,-51</points>
<connection>
<GID>23</GID>
<name>IN_B_2</name></connection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>150,-51,170,-51</points>
<intersection>150 1</intersection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180,-51,180,-45</points>
<connection>
<GID>33</GID>
<name>OUT</name></connection>
<intersection>-51 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>151,-57,151,-51</points>
<connection>
<GID>23</GID>
<name>IN_B_1</name></connection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>151,-51,180,-51</points>
<intersection>151 1</intersection>
<intersection>180 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-51,189,-45</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>-51 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>152,-57,152,-51</points>
<connection>
<GID>23</GID>
<name>IN_B_0</name></connection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>152,-51,189,-51</points>
<intersection>152 1</intersection>
<intersection>189 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>153.5,-92,163.5,-92</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>153.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>153.5,-92.5,153.5,-92</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>-92 1</intersection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-38,66.5,-34.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-34.5,200,-34.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection>
<intersection>76.5 8</intersection>
<intersection>88 9</intersection>
<intersection>99 10</intersection>
<intersection>155 11</intersection>
<intersection>161 14</intersection>
<intersection>171 5</intersection>
<intersection>181 6</intersection>
<intersection>190 7</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>171,-39,171,-34.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>181,-39,181,-34.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>190,-39,190,-34.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>76.5,-38,76.5,-34.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>88,-38,88,-34.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>99,-38,99,-34.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>155,-60,155,-34.5</points>
<connection>
<GID>23</GID>
<name>carry_in</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>161,-39,161,-34.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-25.5,168,-21.5</points>
<connection>
<GID>41</GID>
<name>OUT_3</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>159,-39,159,-25.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>159,-25.5,168,-25.5</points>
<intersection>159 1</intersection>
<intersection>168 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,-39,169,-21.5</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<connection>
<GID>41</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-27.5,170,-21.5</points>
<connection>
<GID>41</GID>
<name>OUT_1</name></connection>
<intersection>-27.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>179,-39,179,-27.5</points>
<connection>
<GID>33</GID>
<name>IN_1</name></connection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>170,-27.5,179,-27.5</points>
<intersection>170 0</intersection>
<intersection>179 1</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-25,171,-21.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>-25 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>188,-39,188,-25</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>171,-25,188,-25</points>
<intersection>171 0</intersection>
<intersection>188 1</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155.5,-15.5,155.5,-14</points>
<intersection>-15.5 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,-15.5,166.5,-15.5</points>
<connection>
<GID>41</GID>
<name>IN_3</name></connection>
<intersection>155.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>145,-14,155.5,-14</points>
<connection>
<GID>42</GID>
<name>OUT_3</name></connection>
<intersection>155.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155.5,-16.5,155.5,-16</points>
<intersection>-16.5 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-16,155.5,-16</points>
<connection>
<GID>42</GID>
<name>OUT_2</name></connection>
<intersection>155.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155.5,-16.5,166.5,-16.5</points>
<connection>
<GID>41</GID>
<name>IN_2</name></connection>
<intersection>155.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155.5,-20,155.5,-18.5</points>
<intersection>-20 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-20,155.5,-20</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>155.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155.5,-18.5,166.5,-18.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>155.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155.5,-18,155.5,-17.5</points>
<intersection>-18 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-18,155.5,-18</points>
<connection>
<GID>42</GID>
<name>OUT_1</name></connection>
<intersection>155.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155.5,-17.5,166.5,-17.5</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>155.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,81.6,-90</PageViewport></page 1>
<page 2>
<PageViewport>0,0,81.6,-90</PageViewport></page 2>
<page 3>
<PageViewport>0,0,81.6,-90</PageViewport></page 3>
<page 4>
<PageViewport>0,0,81.6,-90</PageViewport></page 4>
<page 5>
<PageViewport>0,0,81.6,-90</PageViewport></page 5>
<page 6>
<PageViewport>0,0,81.6,-90</PageViewport></page 6>
<page 7>
<PageViewport>0,0,81.6,-90</PageViewport></page 7>
<page 8>
<PageViewport>0,0,81.6,-90</PageViewport></page 8>
<page 9>
<PageViewport>0,0,81.6,-90</PageViewport></page 9></circuit>